// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ptFyQNV8XfkYiFdANMbgB8qYywUv33WqQksaXoaQuYeObTNeH/hYL+pgFhjrYbjt
Vk5cDyX88XWwj/kHRNjA/tRJyuyBRpKZHigrWd//szGgGGx5QGY3GFDsMmAZroHr
2218otOKF8ddf1QnntYK6a0J02Qv9QnDvfS+dinCa+M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7664)
GFGEiAJnUajVd0SOoJsl77mPU+KprV4QWfoSdB2B70ZMvtgwOuzYT9FVFIn3zPcp
Tqtp/EJByP1LQpIwtdbeoXQGwkhpHRInJPKDO28oRgmQTKxrpJPxdSN8qlh4rVnW
apP7IBf0fjwUfCbME/eSdFV4qu9kVBk7o/ROnDrzUUMnzERz0OE7cMut0XfHW14T
Z6zaXwYS/MhnOs3Y3uFktvMS9xQqm8ykJE6B+80Iq4yHIQERqKub93mxrkfe1x3z
xjTyZHxT4Tu4VDUAgvkKfw70+mZE8Rct/2wmzM6q4coM8qbuiIUBr2Zc/RfzCI+p
3aSobqruyyT776MlrVSBwapCqUtQzKG8VjXfhXNZzeVvaBTiX9zSq+vJs3X0Zw6t
oYDuI824nQej0+q9YGRhbCndICidJQfGTLk03BihAbNTjtdPZ9DuawNFOLIfF3On
Ug+iRNnZsZMLxQR7h66DGgF+Xcs/7cgmv9fgoB3LJFe9XwUfTSQvsNGV9pwwY2o1
WNEChKJc/ki2KZMKXi2z2LQua0dw2kRDS6FyQBI8crPW6EBCWHSdmqQ8cZ2m7isb
C8eJKgihK+M2C7eAJdyuIoz9YZhWjuE41n1G24fLOLoBSzDgpoOqhEFb98qlfbx9
sQRASK2kX79cb/Az5DCSeXTknGPN+WYFR5AkoSbcA2UgUiqwC/AxEUOZ8LmuHay0
PWSFlMuc8wvXt+Diw/njBEX3F3Ug7zyYk1SRZxHEjtxdu/J9UVr7Hyn3EXcFumWk
N47NDT0f4I8nxtiJ7rMCxjACUaBpVGhxpLfOb7Kz+r6h15gx2UPCspATAbTPwHHh
E9YJfK3z28909LTlOHQUylhRtKOK+Lz6ZTeIMq0wnq47mXw8cdXRU4laXUHn0+Dm
hKlOxN4ZuQ2u3zAw1KmApj2DCUabvuckiq1IEBesz4JLq50lzyYsXk5pSzlGccph
S456BYhSEqiHVHKxXUFCA4qQdFsd0Z8H5D5R2IgwQqH65iD+Zw/UgfzxNB/jsuHo
gyBT5tw91kQY9iKV3i1DleTxbMA7obmrNZ2mXsbMiUZ/G/8qFRzOfFiC9BZu7B9n
goOSoi1hB2Gb05Fu/Wgs042CqeCNUNW7lpZHf3JCjkXaxUv2ZLf4yl8GkfGjkrK3
THYCRDfbBt8iAWtqcS6jSzZnmdXN0Bx0D7Aw1hLIMqXCWBMw2nUvFsgWfIOGHV/h
EUYIOW+govj7zGnrl3794gxNi8NYJC206osH97odwV2J5kqosof4epaDdgqaNd9y
sJWRLqMEC/OtomJAPmBYaJJn2St11JDm73Nc0jSXwHOL3gyieyu+naHaZhEfwT5i
0ZJtiT1IIOtpOycUvnxjRCLciHJ8VlEGYBh13DYHBp6k/s9XA39PTrFmMupU2aO2
EKRgp/c9KGyVjgMqasWxtzva55YURg6TEtvdA/L/KNuU2x0y5n5eDSSTSHCXYWgS
/RQj5sE2RHtPX5bbjSUqOiK9qOasxUej6l+L44OJsyo5IgYNWBrKzf84B2qe6kcM
buvp3wk7uAYf5yhjrvfgFw+RGu3fVEbcsps6wmHvelbKmpLSgKvQZld9Y6pJbheL
SGXvlXErV2AIKyAJ3AudTJm3SVhk5w4NpMp/YGx3C4cpwf9a0gBbU6RbW2UHCAFy
l3pwwBKvooUbDwX1A6H8uPwukr0Qh8SpVbJGjsfnGGYIy8rTPF8x48KPNDnqfBi7
PS38qwBVBaeHgPKhCOU94xFSu+K9WNzLbzeB4Yz//g4ledENBOjyJaARpU3yTZ29
8ETftlOVhU6+2snJ4QbPj1JfFurlndqb8X1u/1AaPZ2Timb8zhfyX2GXENR83aAn
DCHlcR+cPjLth31YBluWi7zNx1S3lsiJFNIfbIbBU3cX3S7C34B+oDugIz+YUxqc
6Mr2dwfp62z07qEaGNPatyuKUxXkLlgy+XM3vWLwZRSeZ0h5Kg1T4YJ+OpYkMWNq
snJY0gJQHrGXbv1Uv4EPHEun6Tc7vZ4i9p6hYdeiTNkpkf5R4/rZSt8WiqgSpRqN
3RI0hv6B1oOZSZNb2zHmxCZ3Mwf/NJXMQmV14RINK+DXtZG971DlgGd2R36o7qBz
2R2Q4lmAXnJd7anyAAUwuZ5WxUBygWJuMmo+Kt5QhYZlu7N0mDIN34EGnO4/FBL8
s8a2k7OgCSOfTfYCaT/jnLr2Lav0hHKQXt1pSA+EYaXkuUzHCiGaxKYEHE13mA7J
b8a1JuOEnT2LItCAg0os2oEms5c/0KOkcDxLvmBxLRLGrNFkduKoJdpCekrKFjFM
2lIMbN9lvGnzxCQJeYWCU95XtzPHgM84yjIpEDs0ittAYYyQbeic2PhDlkur6vht
9WG5UpEMl7lYoknJ07lufFNJr5VbE/wRHNHA8c5JUWMtDY9X2PnL5NLzNidmwxvE
ZkSSOVIzuNNDAIe1W6We4oKyoQAHVOdAt7YNx7+1HzqxLcIzouenRLWG6ZgzWHVC
Z5U6E2ueKHwHfkwLF10a+HLPp065DtXvkkfCBrQibeqZMA6sGW5B0DsQj1w5U7Db
2c0fXnxUt8L43Sz30Rau27zE/oBzegThGi4vQ/MHhIp20/MyxjXSNyye9ZrhL7TH
o8hSKRxSfpb/DwQN+lWmBAyioTsAzM59JkNIQ1PTxp3ihSqsqm6YvNmLUuEGXe8P
/XY3s0NlVgvHvkaNRjJBEozDOilnrwfhAp4QAUOFIXRGl7IRkT6MslkgRca5nVmh
ZCKhWff+1+DSAPE5y9j0uOmgAA6NFvLEC0x47zYS+aLkqR2bHGZgbPu7zNJ/ZHLv
W76MilxPE1JV/ag15Nbe8TDVS93fiRMRelcHRM3sOXedkTneleqiocxRQeQU7PU9
WSSb2Ta5HBmTrLJj3vHyVvTP5BCg2VengwmKIqlmFpTiLBf0GM9wrF4IlpPX4sh8
Fo4rZo54xHS6Z6+3Rtgze0PuwrVauupcD2Vmwq8Fbdg/Co+zqQTFVOrOjg22cz4t
N+jc66TV7J5YpPGyPMHPtItEKQRhvvn/4eZSkXSVF5DLY9yZ97vx3tE4uNPldW9S
z8/ep0KEyYafxaGyQV6SYoNjxSwyI+aKPBgKi70T5QMtfLy2fvaETPtkQSlgHE/3
80TdQQHhAAAbTWsA1aL/dSUP98MhmlfZoKyH+Rk5F1/MtqbAGQC2Td0zTrLB09UL
NQhhkOZrjaOi1oGR0aKvzjHxb41P3ySN9K73Sy+QwNA0B536COkJopIKM3EXNUCv
bxQsX/dgMMVfVH3lfdoCCqaItaARiXQ3Yybs5sEn/SptPPJpG25b8JOuZVkO+SeO
6ndEr5zF4mZkpyXHtu6veVUwKfwE2OFfy4gNAQtkGUpcZnRsx7MpD8czHIdDKzg6
67YNsEiaU93bmYbdsHJui3fY8WYs8/PjOLbv8teOgcgrxT7BH9djcB6EcYcr/0m3
61LgqRNQ+CAxctiRElTX0uBJce/Bq3MVuHZgB5++/QpKnK85X5IonmaHM7LRKEzZ
JDdlFLtAF5W8og4gYvg9spOd5P+uFGHNRyil+mMxw7ikNP1J8PN3Ot3x581RHKrD
dwBbGZam+AY4y1s/3DdrnTU/gL1OrHH5bXo37ys8Wwdty/c3LWSOrXxqDHO0M5am
xYjGtDlkFlnIrRK6HEo1J7HzRvPoUOh0DGj1jTcFOMuO3MuTjgdA5ps6es3HFK2h
7s4j5FAhl2mLdEovDewu3J9cJfi6U+5YLoEILeluYEj+Eli2yrHg8S7DP9PkTkiG
qL5pY+0nqrQbzL4g6bv5tXGJrc5EvG5VE80VWDL9D4q/Wy1WHaCXn9iL7BTEdMJi
sbG+nrPheXFE+uuNgCRF3UhX5hZaN4b174KP3wULlQ3Lst6Z0z/ttN3Dl0iV0Jhj
EguhPgVe7dtlV/mW5pOESy4b12TxRHSlnmhmlx73DSRY6wDUW0io7PbAYtW1jLHu
Vm9iTjCN0EL3G34Ho5RmVOD5u1+dxM4nclexFIJN8FTMpmhxYjceWmlMC76pnwsv
cT2NBxqMDM+VEr2+zMmAgRthMbY0Ycsybde1Jaemyexr1e0Evd73dt0ogcN9evXB
A/NJhTXkDpxBYdbULIIg3Kzif0irztfOGmGhO2HeRpfUSVXz7ddT40G0A0b1NZu1
W3oSldAY54KJKiZW/VFw0QS7tgQGocdRkhx4w+HpVFYemeLZkNxPCjBrOfJ2GDKJ
oKNc8j8Z52u4D/9bgfdQKkTn1q+wWESXDnZWtu4h7tF/6XHGTl2FRlE6GCSqyQi8
W6WpHJ8clrbD7YAolP6Fnq6dvP9+9MxaAxuB2Z0X0AXRUotUHTfr+7WCgjloIozQ
/RE2oEjnZKbfladgYYE1gcvSvdsg0l9Oj0nmn6teRSjm0Z23XAsaPkO0V697yeEw
Pyx30uWvk1uEHzZCtprDWnji8nrLjs64VXGyjktym5fj+NA3X159vfFILOgIrDmw
P+lZI0fqiy1C9ngReXo+mVvUckLrbWXlb2fZpuqtta4MArIrPASig6SnNAHmzZtb
H8/MX27aQq2sHQpWlXZtBZpxLgplGu8DmU1WkP9LIFWE7MCKooet1rS9rNelean7
mVxwBTeXWiL7dWJDK5GhKbBhB6lbAcgL/jonXfSRdwCVUL2r+VZCLoPLM+dmEg9H
7cq3xP6kpbc29vgriofF6FXW6wn2YZ1HDW2cJSRWVQQdjXBFMlpLo/u8hNc0WcL5
qy3X0AtZHHXaeMWP8N5pLbh8A7MO0FcNyF79M0tJ85Io9d+0PxZgzJ49yt4QUnIa
dGjszgaCOomWDsRshtBqRoxxcboeztt8xgeXNu4x6BQAb7EJUHNMb6SDO1usNumk
pvG+Vr1HItzLjOOBvHzLD47gwZnvjoaEWwhC8/DugZ06JCXa888NCVLQ70VOtpfe
NbIm1PEVK0p7wwMb/X1exRcb7QRR4LnIBDPyqrgRPq/+z2MYHO2ZXrv9OTl6w9K3
14h8LAqauHaUKsOR+nyZVjOMfer19gqy3oOc0GxF5/5OByEV/XveKVIoM9AmbGFN
ltHTO8W7BkfXypvCO3izy+r6cFDYrOFbr6LfnljJFGpSwHVLe/vDwtYPojYRfRpu
WUJHh5a+k/KvScQ1I1u2/JrZN64SuG5aDM2XMohpZDB4gfkwFx+4gcztc1LXLP1d
uR8RHZ2Y/goNK6gDGRpxgB42FFS+9HYrGla3Tu5XWPJp1RWJ5P8aOad2AtXKH2hU
AOt3zDerAyYvZALGGlqXVBnemqOQpfYF2mU3idGdKkHOJN65IrTvqjOVHYRzJ64F
v4vfyG/ICFR0J8DZnwwDGjywNVAcnuiRthE62wvPKS/t+Cdgqz2Zl3lERDwmn1RV
bYDauFi+2W4gNVhbjSUC7jOXP5bfPJuFqg0NaALvwGQ7Bwlyfnhy6XuuaJ3UE3ld
Zc5qIODfyNNR623RJhXEVcqbIrgyc2j/9Ol7r9320gwh8bcjzalpj34iOrSNn4Ps
edAUqBmg/rpT036/BCj92carCKQc2KLEedlyWP1jT+Mr1clR9uX0dZ267i9KMh9h
gfGhPxc8gmBxvOqor/AfrUDOBTNmFVTGw2uC+9PtmYsPJS9tA9b0qi1d1XsDhzYn
ymTemJ4BXdG2ElNm4wZojDgUgFMkt7sO9lAtWzRwhZ30U48U0aWIv/arvS9oQ5Pj
qFR+6vGEVcApPr3ZzFbZkFfMz6Z0zZQIyilZMBjDJ4vZZQJoORd2nkwjP6uMl2S+
2oW2e2DFpjXiuNavCTwh/AfxYYXMvxIajnm1h+rth5MujThdT+XvGYhIJSeAm11g
8LfZeBucXiMzSQ7rURJXZGfFJvs4e2tni9MMPLXCbmtlxMQZgFsd2aHK7tgbe3aq
nT2/T7In8l2XCX9CxCUtP3PQ6Pmey3G4udCYSeRxY+lcnPoG/dsh+cU8KV9RzcPI
DMKvNMUli3f4JsFcSA9KGIpVMCd2LFHzNiJk7ndJe8HmIk3sNHyJcNWt9KR78UXl
UCNbFOTVYmYcHPVcPTe7XYCRpNeQjMImU4446QjF4UB1pyj26y5UzsZCrSxwHzUD
nixbigxSasYaNnUURWhRASqGNT2QvpHnhBrTAQTlOLN4TTYbRY0Hsz2GhEvzwaLL
wsiS3lYdhC3gu2w1KVGRBsaPqjvD5KyDmbip2nDJnF/306WpYqru/Ycxdev2VFD/
KaiNbI31PwDLKhOGrJ+z2iRRBrysFEgnmKYaz7FQScPyF2iET4pqbdhhvXTWw3k5
MlIWBjWfwGOIWWtW6zhYqYrFH1+QV4ZoCif0TmZZD7BItO97vrLk6safZmEkiaA3
hofB+HtwIUn57BGHjIt8oE3KvplefwJ6iedUpE/qxEYkO/O+Y+FPj8jzr3F7vF1a
Lwtk072mx/x3z5KNPzoVB4UcnSRjm+7tY/ryGLId+DGNqTY0927Jh/8CzN3Hlp01
xiO0o+lbBgvVUmmNll3MO6Q/Noc2hN93I8k1L/prjblIVdykPIfefFZYxOvH8CeL
JuMKlq2uSr1vGgcriDFD9gCJnuAHU7Ap0bPi6xVzDlPcKmmlKZ0UlQH9ZjTY3veH
7cAE22MLGpN5S6NPwi8Ea3ibG31A0L3OcwILIy/NOjd81wvYGCledfsvuFn8/e/s
k+76HnCM0rjGMqfmBZ3+1FmLq4KyOAvItVOTfVwe2+PtfPlf1LpcbYtDAOHzDDE5
VngaZTOqQk8oSUJJPl3WNCStWXdssPpeAcSPpGErPWLBDSPBNeFx4X6ciQlpsgn1
DzABE/bgWFQkNN6wqVuiBGJsqAXF7qyEq/G84/baZxm+t4lfrcBFtdijuENJsqbm
uZhmvp3f4PkJ+z+D4/MixGwQ6dFsRBLs5EuHDjBwLnMILoqz3yiVziU9rbI/ys7y
cJXX+b20wokG4s+N6rwcOHjt9wUODpmu/gCN2fEL5vssk+wUtVcp9W0EScBOpcbt
IkF47gCtLgqJJhV7cKh0izaRAayJlEPvuXEJl5eFos8CZ+GeQ7gOMQgP4g+hELWi
fV7yWAOh9meyjj8EicG6HClB+IEXOYUfBq2NGWoG7EsNU8vZ5EAcWKWfTinJoNNa
z4aqvzWQXxkir63ZrZXT6e24sQr6TzdIP9NprlvUD+VPBfAUjwyYUHimwHvvoYlR
+gZmuluxa+CulZK47RXvxGPWtmjXnt3GLtQ+tYHBuIoc7hgWJNZPxb1mJj76xyPe
2RPHqeIUTM1CLOdDD3KX+HtWgADi9lC6WNg+Hcm7iD7k+6xalZQKhm2oDX0w0aCR
S/jcMAVrA7fICpN1i03xPzptZOuGZIRS7UVmCR3LQEUgj1UepIUoADNKHvY1rORH
OE+SQ7DCuYyg+56dKld0gi50WVP9M7y9nios7iOb15HT3oTBXFA8Ncvy+UBRnLRO
kz0iL/J+Qwbnc+oEmcLmCZIb2+GfPZS24zLyP5ncM0Z88XXH63BF4EV1JFEkXjOB
BCFLmjyhRsZTgkbdq5f1E6ECKbJ1j7w8bPv8PYNCcsGNm/g9Uw7ToFVCizrK90V1
rwHqwmHq8Y6ujbEUPfWTR3hfBdvkHgbB4Q5m3Q76kknm8D1rtvcQm+ErUGd+b0bK
weLfOwrmh8b/+ArmguPKrSTYc0l1pgMWH8hFrMuTBT/vaUrYJozqwtALSlw41srG
qkzZbTxeRN55HyPFJZ9sM3bGpB1ng6/iHPVQI6Xqy1IBZ5l9OchSFlrfWmSG1HCb
oYQtjnnHL27kEFTOFWM525DD6MgPxO5TSPVd0hKCLirP+wmOlXOZujZL9k5NX0WM
gZQMJXnkpCs7kppxSFAV0R6BusLUeshc6pLLL2m1x+OnVWuvRH/EKcLYdsUZs//F
5P3WEGTQaP5DlHAmKnBQ5jakUWY7vJD7o7+3Cs9DWHhvNWwyuwfqGMpzr++N59Hb
J52KldPUhTFZF2zD7SgbWag9iLq0VKmscLEqmQ61VICcmEQrcKwrI6ejr2BK5sfR
fEMNJEHZwQYjyVvINKjJ2shQeNtR9iNaHHCZeexrwVWjwFRjg0ljRrCBb3/8qWVp
DmAbbSsH2cziAgYZfFvhlb8m8fVlk/FRvBkfYzJ/jAr8+jwmIUYMBhi/mqOZlKaN
WorodAC3E3eMykxXZYhMtX/rQUpZQa8muxC+23ERSgN5AxNAB1GEKsM9fMmz6JTt
pRRvs8IlbyacP+VW0BCAPdcz6Ua76ZHjk6oUnzGmANMD34tEHss23QrdNuK+0gQY
TdiwONPE3OyjSBow5hFPEB9EVb+jYh+uwe9/ReYaxLiM8pjve2nuzeDLPWAKvrR/
PkenqjU5WNqQOLs7wjThn1BkHYS6DVnix/J6IZgF/sKslfRlGtzTYqT8Vzwycm6t
zR3mCKI1FuPKMMZG1/zjK/ajl3i/PXqRIW8B/vj/4PpLcBPjC8b7EaQC3iWrOBDx
YDpT6uwldA1FFixTUhQCp4znDCam9AuE5XZuaWGQPKNw85EWq3H34TtdXUGl283z
M3L+Wik/OqtP8co6jlcYIM+QcTxRmPnL9JTystkBMd8v1TqJjPUk9OOnTcHBOhl0
ikuPSOgbyxaY9+qixp7hrWR8+ktAqGKO68SVHbMYjAu1kACnDiEexlG5nolIwaRa
o6T76gmyYInFqSMjX7IPxl9+s9zt/PNIlZw1YHu59gqQrUyJkYoOo94h0uQuSQsB
hZgtGvD1a14HuNSw8aBwaaUYOvMJstUR8Re0Ou+dFhpS6WDU8QEVT6Z1KpjFRHt1
T8bowrUm+k8U0uxcpBzfaJnV10JmW8O/wFG5Qd/6u5Qre4PAjrzZK3PMVDPNlCQU
q5ti7hSuTQJfOsG8tnvCgoFL5VGvg/mVtaoT4HesNhKXEH9V0u9Yyfz+F/Hg2paf
J9MS/uUbf4ZOmBGVY+mVDLQTl1enPbsen7yF80dQgL3CqBlxuHNx+P4219dC8UeX
V0bDhOyDCtDKx6k5+qnUsIHS2N52GwAxP+Kl3k7Ey+IbUi82RjVTwOYQgdf2DsXV
KWH8H53vzTnwLeW9+Ll1AgBpTMDkvH1hDpgy+0eAlCSErVtz4m7Za4xV+Hsgqarb
SfrLDlDW6y6X5yJX6uPl8N3nh7OZzPG17mQYw56f5BcPjWDhC8ol+h2n4F4Mc8HZ
W08OdpbkAPC1lUsFzV0BLahi6lrzZ3NeHUm+nGmPCMAuJT8Riyo0in/5PK+H1TI9
B4WOvB9ACpg1X8h5qgOEL23Uu/OZZY9HrhmibncNwDz2Q0X7dCq+UKX9a1D3PsOP
h+VVFQVb0wU2Z4YWW54FLCX2hsBMbgOpkH7CDDSlROoTy+4ysdP790EciWsQqk22
Rfd8OP3pkrFwHxx87j4+aunygcsOpr4ML6ZVYL5ve64NKD0ehnhK61Wx7j1x63wK
44AYYHrmXg1QYMQzOI3ivVuGpMQGHAsAI5O5wU2ubSrlFxebujrEpw8MLrT9MPMW
0k3R/6yKR6q2cdoHHUSo/mAWdwKnQ32vcITGiaB0rixdl5y/bzegGGmEH78A8cYz
FVJZTbfWtWzoiQxaj6/GwbLYmIbOrTig1+PEhJQxMOeVLL3Q5QmTivTRtMoen49r
ZPRys1dbL6h9SWxKUpZOSe1N7yfZnN0poo1ii1RFOWVQtSIM9WkClwCFCE7xDIn9
gT2S4lrYc7v37Y/6Zc6iwD/5UQ2n4hfNzL2RBcbFpbQxeV2j+56CQpWnHykz2Te2
Bwvbi07BJHou/iEi1XVox8MPy0nf75KKnKOHxMUc/lABiDxeyGkCpU0tG6g15SCV
GCchS5lsiylZbqb0GyGZS26rp3u6Tru5hVLCtdpMyp523wOJArdFX1j7BfiP1aWo
W3fUWKsSQWGxYrUufHJsQkJ3dG/IZwf/TC7LE8wSsLd0RwoFMYHAE1QKy32rjGvy
/cMnGnHUxOuVFa+5KuIONk00pMdi3/sAw9uDjIVBVIZLAWa+1PIM2AfFCtw6XVFH
3Lfi5/h5hSYNaUHsrYKp6cf0vzZz6icENo6zh3z8XsJJYNMpmeL4+G4/yll6SIyM
vO5ewVBA08FdSd20RrdrYN54bkVHJx/DBFmoNMSy2FtU6DwJhA6gGe6j1YWcb98O
GPVQgYAamW3OijZrRvdDkg/zRyKd3ZroKMc4UUFQgFglIyr82l7p1h1PLk62vbPb
QRFeOKVpwMvdVnS6uWdkxjP6dxxVWq47Hk3g8Q6gaV4=
`pragma protect end_protected
