// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MuH2DIaJjegj7ULltpAqbm/sLIc+nIqpJWum33Gmjs0zagj3sVpCl04iKpNwPtWt
Q+jK/BiqzEMzYMSZ0COI4uTR7pS0Gv1T//6rXY29/hoE85OvgrBRXbTkS4VlfqTe
XC/WyW1eA1q6vp8er0Ud0/Rhv0dpkZfKOiPcAwa0cd8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11520)
pzeu8BH7FUItNFwQ0/h20jMlbrT3uEIbTGN2ySmz7irJ+TTr2sJ7OXgN0vZYN77y
5G7agj7JTWyW7dtJOhKw7VuL/OtKqSl9qJueyhSOGHA+p2QA34/j6Pk//eUIQ2o3
qFG5/O4e5L2z89oL+ExcR04gQSNAYEauj1F8lD84MldWGfTReCBTRz58NcT4F33K
GYu0/jiwpTkRO8QclKZnGMe3y3c2KY76zsvbGHHHl7/ChGSKf2AhEb+zN5ZFy3PM
rqCYVJqUtji8QB+D28cPaDJFdQr90JjHNcJ5ejS4/HscefCd8XmfJqj/z6oKPhEu
zkhpsOqZJQGB1qCX0V6Grn1u2+/sOHlwYjJjKwfNk27P7tqSapl7AtY6vE9Lpqo2
z0DudmBY9wnpAHfIA/MIZiMA1lXgYM463irDOcJLBhQGFXVEuw8k6dkU/iPtOCkO
ka9p142QrRvMCeG3PeS6U2MaMJRlujAEZ2UZwo8lwaiqWgS0qFszeC+4NBFCvlqI
kb2kkVJq5m3UECwTdGGKmPFeIQ0zVfSnsDO/uULjw5uGjhRRWhp8RkjM8u9kA0uU
dCixJh91xU9FarJIO7GDyV97kRwryZpFITX92BK73IqLsBOYxIJVaYMJgMGjsrGV
nXhGmNXLLrgDPVdWimO5I0giqm1w3rcBgtIGX2eDThJZFhJSk1kdR9qVx9hGVRjo
TBqV741CukBh9NBIrdwNO2VxErsIEsQeb7wPmToHlxG2E1+0I84lvlh9eCljMqeH
VSXHGAaR8Mtp+I1exe6iScutI74FnH0XbcrdiE88DgSQbV1b/SNKr6ix3xxlf1xm
gSun6l73OssKL+Gsjwj+foEsj4d4FtWs3V4WCB2F8KhibBXTQu4d7zFXPTXSL60q
VZqCBMfwUMi1M8WCNMu20sGOYJRhWUCPLGe4f3+9/isY2LQMDQmc4TBI6FbE+n6l
+a90RsIVlY3aHpwccuwNwITiXJs3n7rblhfhPpWYRSb+cpcqgZe6f+NP/o0sQ1qT
HSBPVuUF3gXsmd2q34xRyRLSftc2RvxTnlAf3GtSIs3Q+zCCZIo+azEFowmvELQe
v9todcWiKiH2Y4Miu+i8af9bN70IFbTyHfbd28bEbhIC616KcgISirnwN+9TbzG8
f8iHg+0XSG6YHmCRUV+NKX/cA1PBKBUlvXpsESboNYzmMUe0Yjm15by647MMfFUc
4OU+FbpqDn4ycj2+QObNllMSn1UD5SsgrDPw9NxXYZQpp7dPjAq2oqRnocI+pI0W
BI5s4H8F3Wexy5hPoQ95P69LdoSgsiVxNpCWW7OnhtlpKWF1KpJBUjID5kru9jnR
C49bSzvoXAV3vXVHq+qO9kAuuX4pQgLnDp/tv01MHRAC4GQ1ZAErg8oS3P39kmRA
1adzSX3tbRFdwZc0Pn+Dn7C3oFX8XaLfuxlIz9Lk/RkNDtCJ53dkScBUUL7muhdQ
LhVIRYGr1ZuAVi3QgBGP3t1g5+82zY/DPK1z2Er+B8n3oRtOa3LY4665osJW+A98
UBsJMVLdtaD99TUx7j7CQi8Mvmeum8IISuhfiesMjc/cPXsmmiRUvtmqwEUlgcx0
R/kWuIfVmPSo/dReA6qB9pfla25SfYZaJMH35ZQ0R+Sn9Comm8eNHkvNcSxka8uj
z/SGfu3FZafyHq3H9HKlwVdAtMoMrbThu6RBDoBSr7kNDKoSHEMScnCyAj7D/Jwd
flbP8JOWtRjHJSaCCYxDTc7NKjrd94wCZPSl1pyeI0YR5zxcbN2ajIxj3xhR8p08
/Ewm+O04xs7fgWvbZIegJCSxq5sUpRCyL2fZU0etXWcrc+fChlVyeo4lLAjjZV9l
065mpl0oUIYAgUi7h45GG0QVzqE7QX6zlmwUvYackAHipBbJVq7x5BQnrS2ezRpn
erMQIlv9gp5zLZBqvmFb9wRrzW9DMuzIOsWLoGRd+KMrCE+S00RQTxWh2qH/My+U
Psm5R/kaEzHLxzZzEwYzhL53QbKq+hZYwWeI6Rfq3ohK33SsnYY/PydIhxZTZWsC
cparMDK9ycRX3oKkpIuY8hFjgqQfe3J6YJ59yknr0XbWN7CyUZye5+/9SGY22s5R
QQ6Br8Hx/LoIjr2FZ3SUeya9Y9hW5UuiuzC6QRJuW/A4R5I2HwyXel24HBA0uYK5
5uF3JI99r6PlHNolq61T3jE287gkTGYV3JzNfk9aGJt4WueQZwBjuorlzK0GAhL/
thhu3ue7f47YTbNGhjTcThxZkHohKDgX4crfn3Tbl195EqVgkjlHrgyC2ocDwHfN
7NcO3bW1ANmNdEG+B9r92SZinito080Wjdvk2Fpg5+MoWFhumR43gIKclZgrrWLq
q7b3E+SCrjq0Ycg3Ps+RkDAW1k26JWQRaZAAfsUNUqF8zwv7FrbcCvvNK78Q9/XR
B7agux2JhClfNEDeQ5jJcYVyrpZJkbCHzukjxX8g5pCPP4glzazwMXw2pdC3Vuil
Mofm9GgCtUU2wsW6ieX6ijev6jSmfuRfXecQLsQ97Gd7g5hujMeg/YyDHjV9R+7k
5F6QbV37fZlHeyGT2+u8t1SuhfO+9Sx5Gx71RoNUDWU36Y3BLseBDipqCybXh8MB
qtQ1KdB/R6x/l3m94KtjQnTeTma+7Xo8MPkOREW9hvmFHdBxkxAuCerWmBzruBWi
nJ2l3/2muvBMUfMnmeMOcfbZPVqnxPo2ksLI8xG3S8sGgrZUjixzjz8MxkfQF2JA
1nL9TPTQ/Axn0kLmiGn58tUJoRdjLmzTmnXJRObodXsr48xILVCL/Et+kfO+0Nv1
qxHCRRe7h7CYla1DRmrQbobqBFy2uY84RbdddI77KiZjBvgcSEQWSYVg2eTecZVs
2bl98l7DHEQzF7YlaGqlTRuxNzswuGZ7owySJRuFBvmdtzPFiO6VelFLHMp5m+3C
84YDIStiA5vd7afa97L9jajYbsafphoF5lK4wi5ISIjFpEIDsNRkkHvigJ6jz0jy
BIgeYwOO4A6T6xkrs+CNa4HkrVECrRulGywkNXEfNGKpP+fKv8GDBXafnza1Oydn
GRYIM3f18i4oI65/6NKZv0N295ALWgmF8MZlU6x8YY1DOMWiuvVYFHkIzkFn2Fn4
lB1jNvcTPZdz938pIY1tl0zSFNzF0h9PzLh3g54Cv69LVNdjnURkZYkdNymNQKSg
FkZGnjbvpSY7X2ZOrWzUBfknpLoH2aG3/Vao7DOkr/ld47pHtTci/PW6gE4ttx0C
cRvlPGl07C47Sn00YxczL+uPpgktJ7rmUMpZbULgmDiKkFb7co0zkGkuq79AiBRc
HhuZ63kGgEYI9VBCEajRFJAS4MW5jcSl5oyYN5DNee/DV5XwSa9lBh0P6J71D9l5
aYUXDWwPEU6pRp/cr7xXsXSRA540bF1d/pXtIMB1dUGdR6jAsuCMyHf8+//ZsI1O
GBopfrhhqEFu1eCmB/2bjXLuE/xrNbBwj12G9X+dQh9Dl/DXYSkW4OW1DPXwLi5i
Vfzv2EaeFFjLY/Zo2DygYmYNdFHemA4bvDogtggixcld+tvPIBwFxuApIfROaGdb
XYP1ADtLi9/m+fyNbrSd/KJ797AhGiezzR1DJ/HPANN4L+y5glJ4Ttl2aNtff1zW
CKbJ85HWdrC5aMpP5j6JOo0VE+P2Fyl03Y/MT+oK8OcTQKWNOAgVKJ4vzck2n+S2
RcDDOEgAMYZwObIbqd7nyxvSe0ZgoGeWMrMyfQtv6dCT4PZvyMH2q+u673GJxsHj
A/WgGT2OfesZTD4nyLAGZCRNqOgmINGsuQ3rb/dTLkZHi2Ej4ukqiGzmeWz2ubzv
7UIPEEXf4KWoCR9etuFVI2mFymG3hdfVc89PYMAdVaPi5qjukyBBj5j5Ln1HJ7fK
cWupMfENPpm12vnqDfN4GRst+dW4kyPs8rWyIJhRBVO2bgQiF21tXjJtmKT6O+4T
T7KvK36EPSgfbxKG+BN9+YxkTE/o/kyLFPhtzndt8nw7Ethad4H5uSHfGR1fIQm1
mda9rZhpRLRckrftao9GIA96gCrFT6IOu/RlLi8YIkaFWtGutuZ/DFaybHGqEFsP
Z0I9LHkPBmGQksfaQ9RFGMB/BFvFkGdTPHbsoGE1QI4iiO9Qb/9UQhhrqJZRakpD
cYjE1EdDoEVoDf4cKKc8vvVY20i9L4lzn57vAz6cftMvbCNpC5Bas6E0wexajCav
/zWWbnIx8UYZ5OV35YRjadakAj/r1Oy5GVH6nijF+PQP13SRd/lBSSk/s2M3y2rM
peL256r/4bj6i77P85i655DJ0RbvX6vfvXc9EoG/zdv3OrTXkNqXii2kYdZC6h6C
t6f1neaaVbEYYIGbsxRbYw9oB1fn9/oTu8uVDRGNLbEthunhrlGOzcR109pL+z/B
fFl5jomOOkUzkZpcSgHyQ/8BITo1Ttdu5ftAyMQzNwpt9ejIv1qWZ9vhpzLGk/6o
ZOKiM41u18no5cWm9cbQcFF5YdkoHvUCBCpuVyXagl9JRNKXgcCgzkf1NPT7/a+R
KB/G1xiW4OQZxSqM9go/867N1o3RyLaLYw0nkX/KSw/csvs6wRa6VpTlQnyZqjK+
VzK+JptRNBX2hcz7HVM2q0cOlVgL+udmjnlXwH9qcTw62aKjY0iePyEVZndAPI1Z
GxYuQiJOCqFxf8lKnSZP5r3rR/QNNqmzdXTKSo+iOxxIv5gYvZ7OoFoE4Imjhxep
atZWH2ykuGgFzaV/uFHX2F/VQVyQwjzaF1S9xFxzAoLLMHJrmVWgmcPriONXD5FP
gJKVPB9x1OR/aMPnP4NgcwP25s63BzMqYT1R+akPUfA2Z/TZ1NW3TpjEXbW09KN6
jCLqiezG6DGotJrQq2gDJNSr6xKS5rE1ZWfXvkjZqk0wzdgM9ozUvwN8MAga9NEo
5uCl95Yllm/ck3E5QIBoTiDNlZvceM1CTui2wl2K+chFJeHIGnyU7xkSLUy9X6vz
Iet8/1UczUgoMIFBi8nSigzj5u2vrTFWnh6qJzZg6qsmwEQ3+TYbwqvAHAHCHwJh
TmZvMHn3vHbsLN3d4nxSyNZVVQEBXYRfGYxMRzadK93ACDdTmp5wo4uugJNAzAYE
udTHYBwWMVdPbZI9y6VhN7J7RO8MB44lFtObCDU7kW4UUJsHyYsAm96U72GuqpOI
wrL8OjPGt/qkmiRVbhwUYS1+KO/9OwzWDPYYwvk0RLB3P6VdkYFv5rHl/sJIZqbr
7MNoCpHZNeOUiSMhw1KsVqmrmhbQdAa7snJhQ3tYqzPJaDc0szMRaXtSe/YebHD+
4cR2YA0sZPlRalSHAbcI0R9DmEKM6ypsBsy6n61r7jWsCM/vkGIleVB2xS/fhARa
Gc5faQ+oKgZ+fiKYXKg1bolMbbRfwMWG+ijalgIUwTr771tohG6Jr8szJn+LJ7dE
xTJMWnDllGmqmAN3VXtuWp4QQcQSuftJwBYXXSI+EAXwnXlAceWA5FPKVmxSreWQ
m8RT9BzsDYlKS/bfwBYZulMFrWpezFhhS1yDLA35FlRTbDLajBlAwS1hgPxq7740
y524XhlOj0kvo1TfgYG1wcRqd71zDR52GyN6wtz/y/rBIu7x/QFnRHRVRqjS8cPB
FezgZ1/DyMNlZO6L2wUw+MEKUBevqHKZMLsv5cZG9SwwVGvyH+wOkR8cHe7q1zxG
SIvmV9Y6cOu1td0loIZnFkGpG4FgvirXwhc2iFRdseUaDx1ooqrDGHa8S6HfTsCv
X77t9FhplnJ0cp+J/LthP+IzoV40ThC1AJCDSoDTc1XP88AH7hWwXHMgJLziDmws
O35yLVPCR9O83Db5w/yQXYE0h7rwVWJi+I1sxddDA/bIRFsYXmlqxxGmTH9l9Qe/
nzLjhmofSwWTH0L2ub7DNai9gldK64d6mO2U+BQcDxNiUxmn2xeIhtwATB0GE86L
SLPaiX9MxJ6sGv8102sHjMv3rKXRNYkVUoVWl3FPLjiQfYRZ70+/oA5dkPwWVK2/
EN3HQyzzKKGX5cz8fNal+2DWXZrp59ZRhMc7J/4rotEqcZWQTqG62ffrCXX5fe9u
2154NGp977giC/kptbqvjl7LQO0iH0Uj9CGARQqF2pAOG7Nc52d3SYF0uYD3Vtsi
slp/OtFf+rPAeAHW7z27HSPD7E/M0oQj1WniAGaKyPKwhqvPWvcHfuVvm0ACdoQX
eYUZ+zFbcQv4cVHBo24AdL1Pp0uj+JD8JMyPZq/5n7h+HAV93IP45N2AO5kIuScm
sB38oKttezDHUDTCmgrEgrwI2a3Tr6vIBYq6fhjdHa2XFAzIJOcswKLLaCfUXSla
VywsJWHNxRinr1vBPoZ5EhjGkqotL0zRbQfdQrk7Pi9XoXNDAMzNVfzNasbr/eRj
/m+a4Q4MnTsVz2i46jYMyE8r4hk3OruGhElu7Si9jgI1lPDmV8u2pnuyDLl5m6QJ
s7kys7FgYcoCMBvsvHFBX93eHR5vWL2bKskPMCcacHCUEu76Xg5f7JOm/tj6LsiY
HS30d9y1viNFfEJs+NByLAnoHQwbGq9s9uPFbv8oVFE/vvY+CyQ4ClP4VQ9qihtT
hLqFr8HOIxF6ukNCwh+da1HygI6pmZbM7b4+idanIc9WFNI64sL8dX0ZQ7+uGRoc
+SVpwGoe4mTcWaOQNix4S7IV6BT43hUMuri0DY3wvVhbOn5eKb+9NaAmFgs1Cq87
nFd7D0YBHglgNnLOrUJZIUQmRC1+oxWr9Dilv3QZIhBaootwDpY4P3IU0O9h2x8l
jorjnDxmm8CI8o8Xew33bONL324iTX9YeJM+J44or7gy7UekRhmQ4pyTttZQ+ZwB
HjeO3Jv+nInjxgLent6a2dPg8m8zNvZ8O16rrDf7EtTvEvbXD9Zm8W0jAVqVfrg5
tS4WItKQeSqH8I+KCi5C4hxBGoLZckKbXzyGwiDvIcVzpMEi0xqlt5X4TpWnez3z
yZKyaqHK5AoS6RJK5rARiyePwI5eEzkEbiLS9VQJeFjJNRWJk0dZ/zqnDQS9XMyF
AZUZB/hx+ZoCPkMzJiSj49XCxhRRRs1Fcwh1I5DRualM68wcz8lkhhQ3CEwS8mqr
ALF68cDDpCHy0F7Sg4qBKc9vA8OlG3qtQtocmygtY3V/E845i+4D0AtGWUiDSByk
LMfNHfFiGnOzdytfJvcibwIZG4BWqGWCbSodQ5gsBaLs2wu5YsnpaoUsxMypLbvp
LJ8fhyDjaJaWdF0U/W5m+iAYWXub2g1sFHVHBr/qED8E6aCTnp3qRcOh10tkoqJ0
Qq2YeoZ4agx7Mz0eu1f85MCdyhsskuLiceBJgIbwwVhVwTF29aa6NTfFqtGWew8A
AI+5pgmz8Pskzmh4V2tgBpUd2mEqcZfs8gK4wENYqkAUSxZWVQs7AZdKSvgyL6mU
0z9+DwME5TfgRST++YpdoGLW1l4iDoSmTfrSfOP10rNcndPyseOoYYmrmlyDlUMp
bIQNbd9J5bfSU8qbEasYSFeX3nAh96KGKtig+8z/KUizQmUP/6149hzxI75EIBe4
u4kPx4nWorN/+4nRa9mk5S1D9njXVKvIx2PDJ3r3DWWsfiasdOq/vcegOAIhHNzs
9zBHlUhzcleV/35pYqagB/N4/6s2Bu6QzqKwLlzlHpQY8BHkR2EQygMrQRFd8RMR
RuBhD1qygM/xaX3rWxKVRD4h7Hzml3D022DIIq3zwfHejATzxi1z7dNTmuqqdzUv
c3Lzm2XjZfEBflTeRqxdWZHdzDLnMSz6YbFFDO7X1135358tp/0v28DYvcYK6o4A
MoyuZ7TPPBijPUc+oOgLrbdQbwCSyNrBGmW//6cF2DrGFl3YjyXouw5sV3gQ19v6
lnovWcGize744AU0RUplVlXDIIPlR8tcCjDvRyIVCm7L/qfzA8wab+1GmK8fEcOx
piJRRGE7yrs6d0ielJwyZoIVUJOw4pyn1N59BzVO+U0JZIhM71s9XxbvN2fJkPN8
7io7f/x7jQGinAQDG1gZtQHVFpKT+yt8yQJwpZPhxMn5XV9Ysq8gTOu60xI3ZHDg
r1Ym9411Nphq9vFA8Q5o/YBwjqH4WBwzNQnfB3i3Twtp3u90E5XIlCzIU063LQTe
L9Hb45wxz/UDQWleW41snmHXw4J1jdfyJTQp05mILpqYIBlGY5qMplhFgS/sPgL8
YgRSpQf9Nw3955Q35sL80UZZBy1Vs0vScmZZptOE1NupNBO6N77yrWkGdQBglhSr
YsGRS9Ue5zyyDdkX+tkOlG8vBP9/dig0VVm1SdYR3xQI2bDEdYPmr4p2jvfIZp1z
HmryGFoJ6BkkQHein49UP/zc7LuXanC4krOvrMkgs9EKGHGILO9z6st+9ZQ0FWgJ
wMPOjp+SkKVvk3gCOQlmUD1x24aegcb3UgEoywg8hrgp88t84xzxuNqEGnHkJ7Iw
8i2NHLaIbu/tpGjDxY5kYjZGDIzoQED+33F9o+2rpEtHz5Oq+P4rU2M8oDVdCuTT
yFWMLGue20EFyQ9HijP1f2rhKj4BfuaVunQH1zFqBM4bfUPaX/xVL+B9oreY9+1t
QtVc3UPt6PLjmeP6jXm/itO4bxQjM8g70u/Lftr3FrYLvAR4e76EDS0pT6Ajbl7b
UuJ+HuJFJtKcn9bNX3PLNXe5X+6uzI6Y9RePHUwl/W/ROMPg9PtjhUtRKvzu91OJ
IYTSawSrjeWxEjU2xz7kvfUJU72UrjqRfTl6Qx/zL8PS5DFpSxAvuvFL6erDcawG
eMs86MgvpXWTvJS/6shzdQXN9988qDwJ3JlCMu6wkhhnAcZ9Tf11LZgbIJhrlzq2
ptU3EltKkJ7bs/PIaCtns9BvMcJz7fgAR0YW+bc9/csQmcqKBILjz4RpjqLgSFzE
A+GC9w++Kkcy+zf1iPQ+eZYpvR17OEyZnKwhaLCb+c7tLHbPoTJxkLXh/Npa1byG
DOlWAa0dLhuQ/LRQxCgxOGFYogB6LfxUZN3JJ96VHOX9IYA6t3IYnedVkQesEWLm
HEBjObr+5KPWrCXjFQu8Vf1N9mUAGToAYJXhoLrRs+j/EXJTVHiRMKIBeQgfKFb0
Qm1FcsfLQftVZMLcZtgmfSIsKHay2nSpYqYSad6UxEfPogkqkkrgjPWmfJNPCAVi
PDtmEV96Ic1cKlpXOS30zOywLX46alxAVnHy6yNzmhE5ZbnHpKj4OVXYdG09obzh
DOMJu8CJ+gkUbDXchrp1kqCRhkOh0rIQ+GPThhBLhoY4vVaynYqcLj8YUbAPQCCt
lY1fRjTAY8gTaFqflWCI8hhtdZKWTMx2o0YD2cXn3kKMbbICYAVYCMAm5JgBWEdf
zBJWZUZoP0Otj4SnFGd+oH5DPYL9N1KgABk6F9EQUAXebGqCwuEUe66l1Tmf8peb
CtAnWY6JKibVf+2E3VnwHVfhPsBzj8dRKzsiW1lzRqtL50BLfEmXTVeYvMcvxePN
n35PKVuu0rszZNv/aYkius36uMArBUQhvZWOvbowWiW1bohQ12S0AbY9lPBiTZGq
XVPizw3W3rOmWvMrC1mwlcFbpbveBWsroCmSEI21lCyQCyatv/1mRodVrysKyxeo
HM2poqZEktsi/B4ZUaJ3AjDarUh9g9ZINWhMNJUMNSK7noBdRclWkc0WBSKmfvKb
+9Rduvc5Q0HA48+uosEWn5whH253G4zy4QK/lS/OOkp/ZITpM2TM8i1zhxFjOl7z
qHXpefNyTn+8kUV3A+vLdQeDqxTHVchITlUqM6seQZIExogUdRWdLmHQDrV2xYhY
pqkH3TW32sDDGGAV6dwQ/YNFOCN7jxYqBzqOB9wgR3L8DlyaU4w3Aa/HF071ds9T
mHOqS77vd7b5gX1dEtbNwJbSOvVtZ70aqzOZO321wlOyX3sc1RLh3aZYpmdKND8o
AkrN20UM8+ctv60Ip4rZmOnovLkk/DpA2L28WrQKAMaZ9MWorc5n2W3LCrb3ADp1
dmhVF8FnKQOTyzkIIDO+bJU4INJvvuX6Q/AdZZEglTL/HIhPYhYFOC4JaUcEfDht
ApLhop3KJ/xJHhVl3rNZnAxayX93RRYm3nkUyITPlJOaDUgXjyxteDURGM2eVEYh
giE9+QkBk5Vyh10s3NV0u1vSf3tSy8SDUfRMJEPQ4Hogy2obtXCNts1bGc6AQrnL
vtufpgJNczx8zZjALNg1knwF3rnTMpfvVnnCFveWV4K+a/5gZfvPevZ/dy86BZLy
44eJX38JaHMNTzqIX/cCfzW0aDNBVf8ID9XBuAbOTKve7Z3mVudpLy32jJJ2hYPo
45svQWM5jVA+c++8vPh7zydTAkg+2GU/O2dAcvYKF+3jSMj51K8wmZkL9KwDtkuO
IdB0lnSnI8uIaZhcUFOFz4trkz9EykuHD+852zNRpAgSlu1zV2TvHUfN0wWTm8rQ
/eedpn+hVBzn4Fl27IQf1KwfocRvTfmqLEJXaVi2xk9ittJTcVKzw/7AtS2pSVuG
X7m8euozH5OgiDqwgPTOsLuTKq62arnqPiUyqNFwpeviOHDJfQrLviHuAiugrl8j
bCyrVComFpOWZKTFhFUGnSblILIe80jW9VccTnuoUPAQ0chh1UE1lGu/flgdq3XV
yLoCWTndwWg+OmrFS5Kg4LoiHWD1SPqGkh1DVVc5LFwKls/nRdaXwOIW5SGl24Sz
wZIcgF9HDrorTFrHq0LM3gTnPARfHEiupX51QFdB1UzMek1N2Xxp+t+LWlzs8MhD
nNwQCubYrZdRSD3V7bOgAWNaHiNOH0b8sOPBjf/qFOuQ0RG1sdHsLKpHNZpQSahY
Jzrwe9Nmuu3c8Sx5rpVyPNP+WT0YfpTL50ClvWyTimkWEIa/hg0dWQeQBOtJKAIq
UQEhQd7l4bK+qBiKNMyOg9Z16qxfT8RiIsExYubLHuqK0ChEJNBZFV7Xjc2msdX7
llOMkqn2bT+o916MUDAkA7gCTJGWk+F9rBOv2p3ZfD+6Jh/8DkeiKbzHen4+sZFz
z1YRq0g24dJQToPeYZ0zmmjyqzH4nLKrXfYP49iH37NmG9yZ/UUExrVhyTpGcJrd
uCky34r6IUbXhO9mLicDnMgGJBy37I6Mqzjtn+Vt4BpvN6riaFrxC83Yuy0E05U9
Aw0y2qmLdKkoHY+1CC8DRPaM8AaL1+pmPfW3kFZwU7k6jjB0jBl/GtnS7weMyBhF
fs+fVD2UoLa7PrKjz5fnVJ6xAH/bfIU6ZmtD8ilKiMnFlO3PGNR7A2HaNU+eFlis
tlAju7SlO0cQceXx1cxaXIkZut/PpW+cXK6VJw2gvfbNGasLSTVp2MfCO6ODul30
Ya0KdIfCaD0cWU83OmqhE4eN3NC3ZOvoVFYYzk0z2a/IGP2FVAKHl4nOM2LLyzSV
BhlmjzQdwCmPAnBESIHwf47RDCtrgQPohypakooYtrYfFpz13Ydgtw098pSYMzEn
pRHfOR36UG4ApGZvbxRSsfP6YVJQYbI9NfNHgScdxnKI3a1imhy1YLwBecX7qFQD
cccJFiSdv960gj4uWTmBS1iA6w1BsQ6DlF4vQ9Ev5Zkdhn6fZWflw7uOcMtHCOUA
R8p6bkqFFG4QYmhX6geBWZMpKXI5sVW6hdLMWqCJJeVxVYpGWghy3ZmuepWHQ31P
TXBwhj2DBnJxDCvQFoYrw5f384Vcxz1xihyzuQ3llxx7Z0aZfxxXRSWBxRukJDGJ
isHFBoQ/rjN5vu+L09cXTUw0ixXlGeGtLN/acIMpaP0PEGfkVvKmwjxIiB+5Lbw2
09XmhWTGBxf/egNchhWzZ1CZnoS+qd8pN1W1wIi5YIPhoOBmGLc/iKnGylm4W4i7
yD7Pj/zqoGsKWLEKSc5UncW+WsaxerBOSysP9paGVLl6QRW1JIRlEttUbsK312+k
cd4Id2LcWP/wtlBLD6WHAfZe86eE+PgbWC4JtutKnZ7yBj+ajP+LuIXFeJlZ7Hpi
6zPDMU6NcZr5lKKBb6yl15+WjezucuLhqBZ0uEQW9WGPD3IzWgFMeZxjZEh/y/gW
cw+wnawJFyAIBPu7GeK/OuFQ1hcrvfJU2GOp0geD+0eOB3dM0mWe0G+AQ1pcd8tj
q+w3EA2EkK73z9y6DJxEeaywVIe8Rx2B6kigxXl+zzSfQHDVJP00ZoLA89K3nCM1
W1aaM6L/C+NyKDr+2XDLRP5pe+nEF6FQDuj6czv3fdiB0vA0PE51bHm46ikteIhS
4zoFdwRTUj40LNjjt3NEHFEXsErXVVRyajVqaIyQe/9YUu5M28/ZWGKzTdSrqbtu
KPdXqkBGKAwGbdfhN0jUGmfbv+SkYPAjkN8fUbNde2WHtp8GxtLhODCn1HTYZv4Q
x7gJ/u6LeMkc9tku65EUtQF/CzrNqkSp2WqQuqppcviVWgvgdp7XBIcMKkdyxrkD
a0wt1A5yajGbE3FPTN7nnidjffzJo2Ek0n1LAZDWYV3nDar3OfZ0WADDtcG15sac
Obzgb+py71iH8YPhdL3+8aZ4x1E54mZ8+OoF4RVELOfa9WMjPkywKGLVSBt0KfN+
sEMHKC6groQgEWY0g1/eCcuyvSzcBddFjMZ6sIhQfiDZNgIMhi3C9/5LLTaHJcsl
KdLEDtKdxrZ8sVd2xcYyrpZsdEvFSDNmF62pQjCLwVfH098aVv4yEV4f4Itq9JVr
md9IsR7N87KzX1ZPcAUizY3bt4XNve2H1UPVQh3N/Ew55ft8yZ+ugYbE0ChRHqbr
Qwdt6uZ4Hcb4lEl5sJhNPIb7ujCn6Gual1MwAXwXvpdVXKvAZ33AX4JRtidK8N7Q
0oB+x3voaeCqdAQTbROqhT8L/cxGjZdnXCtc+4OuSSXpXq9fk340maB2ECE8k32e
xF+Tz9fl26u62GQjPIwEq5/GXqfOby7QowdSnsFJDrqgLfd8kwzhPs75vW1nlqdp
4HP9LY//eQRdoxPpbeaO7ZCLd3cprOTyt8E3CE2bPpoTWCHmYorz/coa3keZPkZJ
4/XJN2cShrTxPyWxk7qjNXZEJL1W/o1+Lf3ws9pAmMXoh+ySze7WDWHR/UMzuLcA
HbX5/7GXTvi6RFGYdBjNlSeWPp7a4c8sxarM85h2JKwC5/2twXOU0sPooA8ej7Va
fXmnr/VufafRkQddCvWJ/RC+Caw253/fOM6OYAJ3M4G3Jz2I7kPisiLSuAPYIIf9
JcygxC/AQoJygjJ8UZgsccM26G3GRBEL2ZVHuj4DTgVjY9pTbC0gcKREBo4L3NJo
RciXZdMpXtzGNpZh6bDxwKSE3FgGMuNrGeqKBaxWMNsIgCfdnunyBLhIPIaEd4e0
lQ79sPVDcZWxxM56o4D5/UUVUBqxwT28LfVrubwgNAZ5LoNb3qkhUPmvgAnLOgwy
ByhOdrUcakVAIlhKYLiof7w6wYzaehsvxdhrs4Ai3nQpMsmSX+zL3fdlNwweAjak
9enaLIu0EMdfgTx3rsrRTT0Jbbxk0YRgLte/xFQhSwa7gS9c3+ccP+U2onpCNPCE
lYTrUXuqYujM2DXyqUrFyGRJyxDCdRlkvPW9EmGoz3LDhPyjcMxIXl2EFoQhecTs
2t3H5dFM57Nbk5jQzTR7as4G0DiVOu42HvH3sA1b6E9zUx/J5za4Ty1l+X3pHqDy
SsYlYMN6o/IG/g7G23GUYtPGWHCez1Y+sQm4MUMAwoBlt6SGplAF0Oqm4jZ0Ay5C
75S+9LnO6l3u6C5C/T+8kkjb6OlrSeOpwtWlYr/A7/if87WAjWegdou1OIxFIE3+
EpokMx32Mz8+Bh8e2PtLPPurUEG4WLAl5nmYGQHA/ezYJ+6oOH3O81Moya7TURB2
BXei6d1IZkkQ1u38BFZ66RB88P8d4pMGUoY+bJyJYOGKZAro4UgW1N6w3GKaA2GF
FW7FHCXBJs7Ggpje6v76hMsX2pPcNINC4n957hYpC9may8SzW1xXb4lmaO0pdoKQ
WlS7VJyvxrtC4KNLWuIFM3/TlSMqpnKhGBvBamLgmktulcK1oQLXLnwj1SVSvapW
+n6pG1j2ZSql0b6xiZA3LCE50tQMl/Lze1lkfqF5igd1mZ+xnrmTXirv8ddtOVYE
M8MwaJ9OjnehfBl9Ez9V/NgBa2rgVEhO3PBFKNTZIe8flJj09OuJ+LKSeAnq4Kql
lWSg0zi5/SurygKdN0i8kYiYaQZe3cYkPkxyYQO+uzMJp7UNCIR2+qoWjnF2ZHTC
8QPKZWc6bevgw0eP3z8p1lWphLRbq5YYvfj5BBDFn6mlrRvaycP33S418dk6hzAR
iAH27mYK52AUkkRaR5bkUEGOuWTcAoQSlSOxelcd9g4uWCW5TqNmkIfYE/Gqt/h9
DEFfI75abrFp+ez+J0RmxtjqpWmbFD0voTLyorxZkV0IPGGOoXR6ROohxAkstFRN
m9wv692HKdUviRYt2CMj2AV05j/O9EIUgWBen6RpOdAdepFIZRQiXa2VyvKt6j7k
nw6TQIyQ568m6mV8Q5s5eCIXToljr7blBRETUlKLhzGYfRXHyDdfct/08LhQJXWD
mb5/vsqhlPbVw3Cz2KrglM7xi0YzE0uFq59Y5bS1XjYxYrZNoGi4vUE+u2Jv1nTr
OO6rsT7JrO+2GR8UQKs6OB6hLw/ceWaH7oqitpxOtArZHlbZyCpJe/kDeQ4Pglw2
6ZZho/PdrEtiRRO31LySAeVNNtvvDJ3XTZqIsB87emCdz6pzfpLPqsUv34LiSzHX
3SdLgr9Ti0pe/sF7V8qha/+tGNTMEM/dT7AlZwGQEe68sSOLVNkhYV4w3Df8LcOd
Yt1TBrOyC/DzBK01NkEJdSrtgaBQJToaBnG3aYhoIt6XdgRaL7myTvWVeZC7u+8u
tHKZd1jA42yb4tCAR08oBPcDgjRC9/BumzpXnSeGZworFK65zgXQ0XAQcm7s0BBL
BBfnLdZNUrABhLGIxDmXpIuF4+7+EvKE+qiCd/rL04SBqXhdJpX+TvwpeUc+NH51
jjJImQs5YmyU870bPyAwiJDg8So/8rw7n702sza/gU2gJBKV3B6elCjXzc5/xuu1
VdkpgN1/Y622Z8G895pzxFO1L9uBmFqSXg/x+UKdj8JUyoBgYVnZJKtPp28QR/XJ
W1UgZHL5RwK6b882BIHpguDpO2SSH2KoZ0n93yCdxK0P8doxfoc4BAcpviO2tpWF
5TM6ol7HkLKiTN32BX8M300JbiCcY5laFP1GotBI8Ax48zCUSJ0SFdG8xvJjcuvd
dm+yv19fP+A/rN8grPF8NoR0QU+n9ZY59v0jx6rMtf7a3+1kV6vQwbq7G0sThTiw
l0c8f4m+8xiiBxCiDQUNuRDrq3SteMj6mjg/2q96FF1nlpFyZINMfRzGxyUX2Y7J
`pragma protect end_protected
