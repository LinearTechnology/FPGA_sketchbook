// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Xi4Va6MPjY0XDe8jwX+4zDHjVUVNlPbW6c5TEIf1xoxpeBcZ1FptaLiccsmvM22X
ADpzM1frtIJ1P5LWZ20MMymw+9nBEx5MQme+6jvpTTRZw0rDyCb8cH3F5lpWP57W
RZHBPS6a8GD4HeeOCQyUF7SDuh10/ik0j4nlNpaqKrw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4992)
+osII5rTdzfZ3tpwfXNzAmDSu/hQ80CDRdkpepInZ168QuyhWBHA8WlD/QKGSWhV
Gmn8WaOtHTUh1vzgR8pERTGuJ0PeTvarT56oe6Xc/ZRvM/RGtnrs/MGJtxYmAMnG
+04VYz8c90lt7Q5D16Cl7dAfEO5t6D7fQQ+vLVtx89SY4DVSlzJ3awFd5f0QL1EX
2fth8RZRnpusCdlo5KVRemtR1DmdJgRGl6BAWfSfEUv2AlMFjaCmsUC32XWI+z7h
OCobDApA33ZbDCIwLBycdZH5SwtRFN2xjSTUKm0EpScmCSmIACWOQP7BUIgTJxJV
SgZEBWpIRVsQ7jUXlI973QZe+czfYrrTY3KDlyayXdGj8C8VIOgMoWcOSShKWXEa
vS9/2zMqj2W6tcaYJWwXVtOcFBMmUHmB7QlHxCVrDaJJz+YWiHCg/p+xIz23lhIR
gyWLxYBggl35XtglyEtI5NZ2t/YyLaDGyeVVFhjV4Pj3Ldk2QfMXQXwSmpPovewC
HgcDfpVk8nB0egq0kl1hHMvXEeJdVxEpx2vEkbHpaI9aXembmSAqB6pPyWnMuFXe
ikhtfOKPqg+F0hdzIuMuOVfx76WwgaGaHfXTAvc78fVMmZgqxfx6Ay2818DiZyj3
QwxL0EhkHO25WxqYl61vpzwKWxi2G7HnE+JbvhYqK9ZaYqt5yEs0B5Uoo1SK/851
zUecS0oPutAzpGQsNIOKIDTTYxrQur49GhfA7SoKNnzotDo8sq9OxM18AHpP8ix0
PFeHcXXTHL1memQYjd0Q8ml8Z9jLo4LyMMbtP6SDD/Rl6uW+gRA2qVI+alXja0Up
iPp6AWzBylnAcezlQCDBHJiWMZdgwbQEatYDVJs1Ky98EKlLYXLcYF0VDHP66W0c
+SJ9zbrmdET8ryY7LFhB0SHXhW4TCH5a2gK5Cpr0iGfm0xqq6hmsKymcWuhM/P8/
jPUbZLpNzJZkZNb9z/XN8ENPNRV2Kl6i1L1eLNBczU7HETFEDe/u1ZNe6UVyAihV
ZWtTIrLuTKljahr1vxyEpX5Lv/hoR1ZyVDCEN3cQYhsevwTL4Y3Cd7MKcg9JX7DI
efpbyM1dpBGpnhA7+NFDddZHooiruljhr7sb1aGoijf09e4pXS65xd/huhMJQiRL
+vH9T9KYTww2As0oJtFpVB3PjP0FVamTXpEi893i9rvFIsYuZV67awTe3CTM59bO
eJkfiInR/HSIiqPwkgY+GuXJ9TBqiyPVZwwtqrjWhgtILcNrpt2gs9jQMefm90cQ
lBdZb2x4YId4aAUxeYDarWoSQIjkney8m7LW+PjBts71MJix3uFtZhcmdWZZe2zh
RW48HgO5f9xVB3fYWnl+vbLEdrMDJlzaqz9YDjooX17vF80n1wNTRIAuumevhlK/
tn4JD1EPnLvghAMIlZxoqFuOgvf78CPG5sU9up/jtXdBTBGgo4ysw/VUR+yo+Oot
yUepZwfywtbT+J6gDKsj8Pt4Rjx62gHRQuLxxv6uhF1iqVVezpyX32mUOH2saC9c
8K046pM2IwdtgWz/e0n5T6j5we3Gy984uEUUFSbOCm/so1escYzB8g43UBOkLR2o
o7PKokN0v5PZh9KSbaQsV4UmSpAIS1wbSfvdcQztf6TwElMRFacTkVYEqIUw4siq
qT3fbohMOnUd9cbNsZfMqZwZDXTq7louyWraa4CEbq23+zwn1UqBE6tGQ+cxKPQc
qZzSa3kFYD0afsW1wLCHVeZ3Jo3NtK7MbCyY5s3N/VoKpjHkeRKg0Sz5en0Mj2RM
kOts3EQXeFnLSWaCfraNbuwP5qogOyFUkkXonzFXp19vJCR4FeVyAdEGNhg4fK6x
GDNdq9ZhdDTnxd3UJB2Adeq8e1OrUXNEnNrBaEwjn3y3r//9gp79hO13azofPCuN
yMMrAVuwIiSZRCmYvhKe0Fqa88azbwKQgsCL+63vtogZ/FkRuxLYpiFzsw5hKy8I
paZsv//IBSbsxOByJk6WgaGzvKmQAGUdQrtX81BcLOfZ/W4n2sRwwmuRNUdlWWQV
D5xEhSXhgEGnAiOHUFCdrQhXWbtCKtzKzTJCo5XJRAla3k3l09/HQgH0TnsO5K5j
DpVLR156KoUqn0TAtWBfrfcNjBzf7d6PuwmJjndVVyQjG3LTc6y34+FKTGOkEaun
wpVVRkq9g9RrEaI66UiV8xSNuI1M9gWMiBC1N8Fv8sqFpYk5JA2CMvullNfwRzCA
Pvx7QUuUiIX20UR/F8nL0eW16QB/Z9ZtH1q3sBCk6efy6JUb/IsZo51lsVcgNMAp
gJ+QX51yS4Sz1bCWteblSpdcPZPnKR6OuXtxS+YyDbCt8bDSe0kZdqicHnP1cyUu
lubUZW0UO+K4qy6M4STqKpFH9bD6H+MwTfvpXTf5Ut/xN48b5H3+UrvuWHcVL3d9
YgNySU7U9jCFOQlz9nNQM8nPSfKhkN+EXa5fdMptPxV1EISNESlsd85nP6+Rr/33
72+TZJxATS70wCMbGVXOo8cxdCAGqy8y+ORZPEEalFhsot4BWlSeaC9kXgNeQPUQ
CdcaG9OL5wuNpa+jPTWSfzD7+eqWmy324F56MZ/O8SJRbEBOjsrEvU70T5YsA9I0
z9dl9F3T544Z8qpcb3sW2tHfRN7fymftbeJuNvfHZrkbWadeuWUx+Hr5dALgLeWL
bodvdOtsO2nU+iuCmZJxOuC694ORMz5l1830vkONvgXj6xXqHKG3a89PiaYnc/Eb
F5DSs5S082m2G2g86onXahQWTasSaMUEQNEvQfv6EZsVl+gb2jL2qjHX6sQm8QiN
f+34K7Z+76idLuU2OXw85MmJSLzGYlUZNKqrdx+cSC8CsgcoxNZdAtDs+83AVdsO
TvyjjGqcL1GJi4th+sWIjamz4RmmJxg2/+f9jd0SS5f9BwmmjR2W1Q5MHizbsyM6
kfrArIhMcssG0FDwIpOGG/cs8LBl17BaawdIrqCW0SfEjn9NMZez7+AkFgj/izRE
vfkBRxETl8MfZM5AC5V5KQ0QZNdd6dEy25gNNVgEoKsf7K6M70NizSWap76BmBKZ
ITobxVDEse37HiJ7YpRlASr4vGs2QVqwuCMzE4rWgnX00G5h4oa7GBilQonk6RSW
GKL++aOTpuI6kHvfVKBm6O+N0lvwcoOewWICDTkRR4QWjhcQOToQXAc/0SaNtlhA
VeJPJw4AmNEpIc5R2XKluLbpMrp3i13WJTQg4/xgaUG/Bwg4c8Zl9/sYFKFXz9NC
ItBdcGiDePY31W8AaLaeP4iJj08cdpbpc26hS7bGzzCv3r0RbVjFTV09b+NS12d1
emKcSlqYBfDPSu9/OKQXPy8yetZL5PgasyIq000FUhK7f7UkjSD2+XsX0Vaosmd2
BBr4x1nfvXl61frDxaTnCA6n47KZqqOUEDtO/zWmqQNtR0nOT3GWWCPXlxoq1LDM
M3MDrZ7IOTzmEBdV+hH982zRtDhKbgVirf4rI4nmlDJRG8857gv+dAMPRLWkMegH
4hd6q0dYDD26uRAFVLxCiBTUiEYtE2hqqwwsap3aZBMmPUO4GHrkuDEspWYaSnuo
bDqstXNMw6+cG8rcWX+Zgo9PBp1iNXF4JHigEFUamaUUaHpoj8pqmjIEFN3qX2MF
v1dsAPfibOqwe5uk93/3DqTqwaf7rFgRRG13hn/QVbqp0sXXAAFCy8d3pFwhKwn7
2b1OOYTXFNmBeplmd7NK6+HuCFUS0xEAr8bQNdD1SrkX/oGEl47PdYztB4nfqh17
XdKj5Y+f1QxysJOGUK+ywoF5m5XYJXskSwwFphylQNyfSjS0T17xFlGILne3pHeK
mazVOuF0O+47JII5QOjB2RdCvy1sbiuGjPXXul4+ifUOxZCMnWbhEQ+AI0pD+2Ic
16QvHXtaKGo6yjVbg7JACxdo7NSnnpXkVVqrrPZ6b5tzBnEcn53iaAXW6RESvTyw
ruU/cOsm+NLajfGInc0HYN4fXtq7WukPtuggNQbf1ZHAZ+erSCGUlhszDb/R8fi1
E2Vv485f/DTWpC7PZ0IyhA54yVDVNjj6z9h8TDAGgGtlRDIFqAzXXhRoyxQs5yjt
VOx258lgZJ6WYIOKal0MJ8WpP864rlfG27UUp1XPDWd15EeV5RCzPj5X/m6qBbkj
NoPrFctf/suzhBoVwazCR5zmJdHkI5UZyF8O1CsXr4uW2iMs0T9NpaZupXTdkXXV
qJmiPTl95fQdZlXKWNhZ7qXyPY2fn9Kn0mXMPcfx2qZb3FUf9uJPyDoht/2r/slv
KqyMuW87REMKGnk2excNAQJ4NZ/iN4DH/L8viAfUnr+nG/Yz2OTor0UPMjfNP3xw
9jn/7ulwXEBW/5wjE4kGM2JxM0n8JAyxKwWB1vmzpfelvtSqySv9KEBwI0m1c77D
asA7+ZUNGqy/up58upz80aCYRMw2SJPpHKjXZwvqZZ3wW9Wbr8uklGuYmhorMsKC
fXeTvE0cRnkdwJlDYMt2m2mdM2KXjuukk6uyL65lPhBElLRTwMhgJENv5/nVjkkR
+sizaad+4Gj4vCMIqcu8wGvgpKy70TX5cyX1SaZQ8RRId687cc7P8hIwHzHYfXhZ
H1LRSmQRWVrDJ5fxAJIILlDuR0WNmq6WzGgSTSG/Bd9FwkarD1VgEV23XtH2hVjP
hoOnsKU8r4MwE8PIZHQcLQe6k+eyEUDRzDjYgHHx33b9y0JwkpLojqeSfu3fOUSA
IsH56nDCIA4xCxhy8FNDjtitWjyRkQtq/NnJpsB2OOGXoNgYepSPNt0CnlGhjVh1
n81oAGoDi7HPAF6rU9Gx+wn7rkTojp0TLZ0Q5UWh5abV9Mq0kMxZ2UtO6tIctaU5
P+6PWsy28NywJi6ZKDqI3RMotVe4G2EfEvVek/x8I6n8kd7MPsiqlJXXdYuImdfa
4xvq7/88aOyC/h4ZqzYcKgczKTdPsng9rNab9Ag01rDegZML3A3jqsfjcjScXkgZ
XLbuEgSbNG4YaW8IxE6BTHhG23VKKMHDVqVcfnlnKL6sGRGtnKLxUfLLD4zVo6N7
G6C5yfho5rWDpr5aF5+Nn8EyC0oXVnotr9to9kQ3yH1YiQypesJgCuJ+m28PMLae
cuwYzmavEDzjFeE6kpoM2JRj4jEMW7ZiusY46F1LZU+6MYvf8b1SdST6NCbY6Bzi
WSPrD34odBxXYGGixhVM0c9LhUDsCdbwKKECW/0l/PihcOvFJQCOmZTc1I01gVfv
mm02+rC9QWqOLYaF403nTz+6OFRJz1BXIi1HfZ2SIHC6ZJ8WQFy8dGzL+nKyaKv/
KLekOptU9oG3bdAj6Scuf+jdRfOiUj28XwU/LbiGfKNCvG+xHKsJnxPJtR0AR+45
t16wvxhBFwQnJqZNvbWC4WYXV/KKXdrxYAJxFPEVXF+tsc6DqncSzN90cGa5uDce
IozOZ5Pa8STZGvLyAjrHd5xGNpcjzN68TtxzYLsadZbJsScGCFUYHKvAYrwSwmxM
Ch2PmTHs2zVGszfy+F3MOA8g0xPGk6u4JihxfNrL0AfU+FA0SB9Faf0bnrKnjatp
+Lm7zpel4UraHm9qxj+vLg7dD+ekFKiwy4Cgd5AVQx+b3c0oZMjFBsfsMpj1JrGq
RYcS2M1HcFlgcu8gkIqRUsP+7/GNZxp2IgzYpd1mITZwtOAmrKJEiXOR24TN/IGF
2T6Qq5vzqRO6O9ji6Iv/LjBCaVGwi03OYTagSsY8mnBZn+9E+yQ53dNNTLilBeQ0
NuGzsRrpv6qn9kAcUtoatXk42u6vRCRROT11IPGEMtw0LFx2OJgKnDtSeDLFVhE1
aMrQOKp/KaC3lPXXKbhHhMx6BLSY4LTD0WO0k1X5dbS1LrzcEEG4Zo9YHj7K/HkC
Vq8yd5j1rS6Tj8eUChfVQ4S+Asxbu+VsoUaj9cwPga44oU8VwZlRxZEHcmxgq9/K
Qe1rrd1iUnuu3NEYafxiIHOAR0bygwADNFSmtZT8aPn+aNDRNGqHQLRhiIWD8hRC
rznUbXqmP3dHhTqT8pengpItS3Nw4U8tZuGCQnqa1D/VJ0g5IYO9CGwwMqCBaH3+
O4lDbSv/fzCL1cKCjnotTP+3qrpv+BMwADy1cYqM0nV+0Cd8VS/SWaxbeSZwoN43
pMbMYxwmf+NZiVNyQuq8uOU7PVlIDnrltjz+36+Xz7sYhalg3GqKfH8BkvXEMjwV
JxJBc2yfKzRJPzepGGxkOIdZ/dZWPH16LpgDsI7JxMzYgSUxvPXj7zeE67eJxhTd
+aaSxWIxuHJU4QXSUjCvfl2IPjAftQaN8v9Ip4qUJW9kpRBqEBjfPmTvUsj8DBA5
MjBS2XeJgxFN164VU4U2icdmKphER5Chlv5ZKgVcWSEkGtXNZARRcVw/7XBkZJHG
S3BN26mK6qPsrrenI8Oxzp0OiZbpo6jkSYWfOa33hrdzHvZKwCYLTBUIaAdDFP7g
sYbQBKCdAeYnt7ZNk6XxhfQGxUvJejUpEIKOwUYejM4/vYN7j9H53Bg9wZ+ixVXu
rPieR3UGd6rV7d/LU4UVLNzEX34MxBQVAcBLfa8wG9Dxv6lVcKtro30W2XWh/WEu
8rQ1JxA4r9cl8198iuCVKNv1lmGTEM0H2EuyTm4hG3CsLrt7foK8TEMropfbP/kL
`pragma protect end_protected
