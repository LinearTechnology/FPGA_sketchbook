// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RJyHAizUFs2zOFiZipC/JwBWEIe/XI31efBLaijiKivFw64fXwxf+uL9yPEId6Zb
yzge5s+Wg4NVwFWxWvA0rQ0S3d1YAiR4aqJ6z8p7qzsyOWz/+qlrItRAyOKqQKtd
gwfua6LSUtcShgbfpLh8b8OOFdginz5GLPPbNkqLdmA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19744)
qNzPH9k25oqCOPly304HP7JmrjsZN6hzTbUTHzo4juocf0hANA2hn9MrPqfO+lSd
WWaXCv2KaP41vJ0anKltTu+nZGTb8FAGy+LQW+CknIuGH2NsKc2xhl8kIZ3U/9dp
dPSqYEdHWMC2gCbzOzF2nTjsD4KB44q2HEeBLvE9XvgtUr9ya3+Hx3ffHWvOwwyG
Zizqw8Nuf2MES/ihPj+xJVOa1xVbRpFB9+0EgC8Q4frSS13Hzn1hvH7yAQF4lKpD
qupnXeEUSFU/ywty1U2w9CkjmCNJbJXEVS9YEzi0qy5szHMp6jC0BsRcDEnBrKn9
gs/9QpSniEbUeRpd0f9qPGWH0t1C7hxohJMpqAkBeTZZAiQnbpnzTK497i5Yf/hM
wFhk0VF9CzmDxmAc4Eh3JLp0/vufU0uYWnP1Duqjj7ZA6YieKO96duoXwTTg76oF
sFtbjjVhH0ZNKCyzYvzOciyMl7OK8ZaIvlGfIqYvZfTtPEsh9M9yqmBSuG8WxK/2
zQq/d+EbadrK6t82uy19fwcL9OFbmeXOc9v70tug7DRKb7mgEpn67y2CFVxEAixb
ykDU3D2EM2ljKFGOi7VzBfccr1DfykGV7dd0EBgGirPtz+Rs4v/Ynz73zoFP2fEB
1enfToR+7grp8XTmivoqCrgNnqZvwWYjpmzBdX6Dnxf+hqAHSj6nBYv5+LdZmdFW
Wlc/oMN6gV8f+dggF7NIgSDZ9AgyiTquXG5/d8V9iGfRzS/QXJpAqzSPQJJ4dZZE
8dSWWDFyM32STQdo1x5w+h2Gdb9fow7MLRytLxvKd/856hfQ/ubN4Qcc1ULD8y9c
7IAWaERVOHTN5RQj37PFiPZXbPEMt2/uoI2HeY01WiMfcKSIbjsw8sWj3C4a6Dl/
1PRHEaquk6Tp0xi5lUCyluetNTPrgacWHpT/fkV2ALgN8ngCvwv54f+AKR7pmrhL
t17hCiG9mYPTwoxi5ZjMfNBRZ+M0izCA3PdkA2rxDD1f91CmmBW2/6ALgk7yjTBc
zl0v4peCSN03xdt9NAMTzQHOJs1q2RyihSCzGkh1MipUK9NQXvbhZCcY7qQd5Qsy
SuaGZjahP2ugUPlK/Vc5AxmX5iwviJKieLvDSuXaz5khqIGNiWd5HZPqEZzryA65
tBVUvodpOyn6wgmPBrF7Co4tIt94WWg8VV6cSneHV1ZZGBrHUqTlI/8p3QbRgoAp
uQ1gB54b+/dKmv0nfcQfVP2X68XKYB5b3zcS6T5DYHh5vm9+sbvzJ5MI/GVIZBER
U4mOrjDKuTanMnw533WJEzY/weW+PRzO3x8Wp+bRwhISqX+WXgh0hPCY30psYJFk
yz0pOmjlKydtoBygithbSg3fWUclk94IfoaPmSa9tkZe7fGKkSnpoc/IjHZJH+NC
HIz2i8y0zWoC+Y3Sr5vM6xNZ9jd+Uvojz/wPnJLyKcbSbzY86tNh1c7voZto9CB3
HlIy7yMoaQgvPtbUK9frU5R5nW2CLyYTuXK1ugWCBxXH8nOQn/sm4MuVeyjDHBY2
ilIuwAjCPNw+P+rVZtt0xSNf3uJd60idV17VBoGtBedsIocNYjIaFDU5gI/kc1+T
EK9zll5q7ndIHU4Wc92IFDQZ/OWo4xK/XCfSC9RGfg3bMbiXGhd0M/Jfw1OgqLUw
/0dxm2ljrfYQt3J+lt8DztjqhjIMZ+k5e2Cp/7hk/PJnJj2cjTgv4Kb/JzPPQF8K
ZGi7pXGLdsz8Hs9rf4CM5nhEGSuHywvliZZIcRGuVh/uhb78JUJvJsIPVxvi04RF
HD8jOjDd3/bnttcdineAUNC/FSTfRHxcAW27iQEvA8cZa3/nPQxif35dD26pT6fp
SrOEY42IRRZcRTO5VJ8lzGWQLl6ijoS5pk/VqHPGNpazAJRzbm87ZOP7oVsxMoMk
cjXHVThZq7p3YsX1+EOvIuThduo1UoC9Eud3Y4YBSpuk+VbmfqtWQHvjMuk6oBqN
vL63clB+H0RYpHcbpq+oQ/uECbPadVjj03xeLdE5cfgAf+rMytWUOw74YCd2IA8Q
gtnwbwRRqQC9ZlLWv6rfHflSZHhRFiVyhkbzHMgi3JRcaSnvpIIzjusdjART1K9Y
UY4/8/tYJFlw/A/lfsNEhOP69fo0Rpi23cGLAkJpl4tBzKv/FiFM5JWUi87P38eL
2SB8WvqlEQtwcZ0OXaur32hPxHNfwXb3U4Ar9nJ1ZwA+Vf5YmMkzIdWuZaGkjnzP
xT3ZNg42IlAID8vt4E5C6rTMpP7IvA/xG0/6vs1PGXQGFB8yP8fY5KFhMTq6fdC0
ixkcoLzs8P2SE0MGTxGi0CXr0jx2M4vILP9DH0zyZX/y2SQ9pV4CdgtyMfY3Sjvs
sP9K9OzaraAsIr8OYUt0YjaYq7Ci0N1Fzn6aC7n/nMbnFpPl5NvWkLixrlpD3p0G
TsVrqraP3MYgo2xxhyX0fdbCChsLAnxNT6teOfhhegjkPa2CXdCYMkkF4XSeT8Ij
demmuBVeA0KBJcyEvnec7wKugZngya3ya2dyAtuBbu6aVbk5MnxRyOi2W3y3wGfl
huJbtefRcXV95fh1zFAXZ0FP1L70VDQAIhlgJiCELVWRMmJwcG2SgtVayQuUV8+l
S6fDJR043A1d9gKnMZlTd5hyJb5ClvL7vpVjoHvEbevInb1au8CwdLsdU7ZN8bVm
aoeWs50Ya1jzG6F/jlB64u4lAEjt4jEB+V639PWUkZtPyAmhD8iOwED09Js84NtQ
qPVA3/wuL2hf2Qj3waCHyryG5ApPM2D1jZpp+2vvn4teAmWi6T0ULP67U+doA2q1
mr7MYvvJ091Yb21eR2fGzc3qs1i8aKBAPk9flOac9gyIFFnQ3bcrVfKt+ulnMc14
6SmVeemqWaeiXTG8/cnyq5RNHUNlyGcI0NThkswu/UzxLPacuuxUE0mYjCSh6zhf
0/IWdAwXZh/R0R1V9jjddHw99E+4JW0Z/LC8UOto+laJuoTmkro1pDyc+v4xd3Kl
GPDHTO00837NCH/7zH+vrWmmbV9vE9Ls+XRI7UlOEey44SucGEpZmOPNEDWTlpmN
7zskzkHAIW89PZK1G+NnDl8AWdx5QPabU6VOr1rvgnITpL505SUVrSiJSPiZezLm
bFx+tAQ8Yi3hgWMRbz0aXwFj4pVRmp1W/d982Rsjcg0LKOgX5weTQE/91RKGoam0
jVRkSBA98S3OpQVYv5/7SYHh0tusi+JRg6XoRItPOamAcZabXebq8+Iq5Q8Sec2V
1VAlIhsPS1eGlwifyEdZ4tbIUpejqB8NyXaW/mnipmqiLAuqqDw/1XcqfedpbSvK
QtsquMC+ZbVp3xUtlPfxRkHbG3fjDX5dnaOEARdHx9+ImcstDI1Rg7+/zZd/0+83
VILhlYyla5NQGTeKduUS6Dui4srebIZej69RupUJHCHZq5JlJYo+e/YUc5XQOBeR
rWKYyXhbmNm9AhP0zz25zBojOqJbsw6skTCbHBUjsXn50fSWPvtAXKwDkMo7Mnlz
dS8ThzF2d8jLh0MI24TV+1BHmYb6cu1w4YMiVgfPBpUIPj5SP/yGDMvvrXCM6+cC
xp2kgvqlsg1y+LKGQUrEfmbcaMu9IAPg4BpHsRGue7fxB1ipGFE6Fx7cTG9Hh+8h
V/cLhcSqzhQZbptecXX6+U5NhwZpy+WuxfQMwY3IPUDrYsiBhRmKj9b7YXnXNkUO
kyquiAPQZ4xuG/nkYENddi+nXZze+ENH/aGpX6zMO2nV4AiXCrzTTiiJI2zlQdL5
TgUnqqq0H6VqeJpdsr5bNtz+dppxMPwwcw8MtE0+O6fn1A3R3C4lnGYdsWqxL/tB
u21b5+vKzPHh45TpGb7iteBB1umdAlWfOD9tt65l4yXaVcC9T276921brp+Y+R1o
b/bLV53F7C005+Rzf3OillNw3OpJxMDtd2NR/gASIkXCdPraKE1aq/t87D/TxPV/
a1G9bVJ4iz2moKLildovFenQ9WQkM9FYoTqEFaTxgHXpRQmVl9q2ZAOcLicpBjGB
Z1ui1ITeH3sFRUihVy4Flyrc/tpwAC+XYrZrBmmWx/e1e1gGd95QOKJeE4nCx4UM
2txCH4+dS4YiUE8rLm09MeHtNZ3+3A6CERkExq6cCEQPV4HdO06T/vOOA0Z6dNIe
qoUb7/RIvz/iMgWfSBkb3q7ML0WTGUF19IvJ2GkGr4VPl4bD3gWXi7E6pv1pWaSM
vvGCvMQf9+no1SZdmYFlxCMixUZC9qhYrEdB9Ksz/zBeREdgamNWMWXTcIofh3e+
oeDikjLj3nDxOU1+tRJ80owTAnHLfGnHRA0M1uUBGI5Slj9o+DooxBKH0YOwdyFo
v0IqKRfr5DzcK94PUbSfhXbnlIsqKAXF3Fcm6CEWLtPnJKrFYrDCzS96UBI8Dj98
Ei2QDmrIrutiCkl0zn0YoaLJEhC03DX4h0jbTtinry4x6+DlEhQ8eW+GL1dKRrsX
2eYWf0Qj3C/eW5aPuYamfw28OmHCSa2AWEps9ncds/Qmt7zUNUXA9SuuYfgaFUay
hjwQS7ANvv6+rc/I5FQJuhAxqbO1RMj3Kvu7D+y06IoGvWZViZ9iy027fO7wXaKV
f1s1zo1oErC/8EziSdbQODm4yxa4QjTPZo6CLC8ErdLsW2Z6BRr1MykDQvEPMO7y
bsLR/nxc6m05MW2KT8QUlxq7/YnLt8xQqVqFw2zmEoUpDkrds7DlRPnR78sQPXE5
8N770FOXYDOOiYCZbEHqvpTPBJYzo9WZgErFt4jhJY5l7sODhWYd15h+it1ScmLh
fWYQTHmxEgUAt/hbGif2hbJDVBJbCkAvkXmu38BQa+B+jfWos0Gq2PAuFO0zYJtF
bhYf5lp2GsUgWcjr+0j7dHD1V7xIxeMFE/zNQ6n0SDQd45Q76UTj2eK20LsrniLx
ehk1LpObpNoBRZgq3UAD6BohpF2jOO3FBADMsIqd97xspL3RDpjblAI7rEPbaGE1
hMENNI7KLiBFG/BpkRzuAuhqNdJE73csU4XdAd8R9OjSuzgCFbtrj0abNsrqd4gD
kB4rnBOHTnqo2M2ZB8sjdSgd85f8nRwIlmpM+GMt480ylWgZz+S+7a+OFReQAqbp
zLJeH+Qm0jDJ11ohKBpNSlgsHxSD7xrKaEK7WPRF4KoZJaA7Fi9NF5Jj8F+2Ty07
mLlclWWE6u3cBaDJ9UCKg7NC1Gq2XNzdYg4fk6UTE58Jl2nyygxYBUtvZ4zzgHph
pp6r/+0rdezeVWkGVtzndqitHI86p5h76jLgXn2rOYeo98A2juRfAFb0BhDuY791
aT/F1xe6/+WlKUu4JUTEEgwh90xTaU7dPpNKg+dAcCpZl8TjyDvdPQQ/DqaFUFl8
OYLC2Yykx210gX5o6xzXVKX8JqbuRB0Q/zCiEXfzZjxnQYfLiwaV+a6XqrrVss/a
fNnLVGQy1c8UtQgyqOTt2OfqnSihpU0VROKXUApFFIIqu9fcUGi/zIrR0zAwBQxe
q1ObFzkZOdKSC38geZYU0PZQTb99MMeJeQvgxee2uGnIB36ri6F8v5pmj11hzcEd
0OCuM9V/6wXZaJ+aMRzyx+fuTIGCsxk/acdMVaGKRVIYOcQU95P+P0j2OUAxJ6DJ
E3+H3WhJH9Rykh/yCNkv2W8B1/3QWZfrlo9+h5WzLudTg9epS/zBNb4uwoqfkmez
tAOCuWFzS8Qbk0qK1CGalFl/ELE4Fb8qlLvpIVRHjKlVyRicQL7bx6W2P9Tn3n0z
EPvb7D150lIcNwdwvBX6DeGb0/DtCmasIeszmTJ8OmqvkcMOHnqdD50uCucqFUDO
nQV6xJ9nw2OJFMhI0zmQGx/rdpPv+s8I90IhCnKGboEvxhQai7YZ+uRIeflhwYRa
L1rnhrmTQCrkvaDueEURJk7r7+QaAiy2O6y6UPSfFtyDsb78F/mRQN9n/2NBcRYM
r0T962h9FxfPuhSayG2ohFBhZGBVKdi1fM9gwUHle7D/y2LuCWGTyWInrb6hxRBN
o1GG+BWK0K1KQiddz96L4WtmUhnywJwYp+oescxPo0rJpbFTebaqfmWPHFvpE8+D
2RxgfAeY9wQLX05sdVBSLZpSJSzI4QAbzKy52KzcGvdxW6Dmqnv/AyfdGEauxOZG
YmDKJ6gA4wswdwsruuMonLgxIFAwub3zT+TnVTb0dxzjMOPHAPT8NxRDO0MvPIHR
E0506qqyjlCEutz6KXuJjcFdMQIhvJrUogZhDwKKnQ9Ig+jqiEXkA99qerebwMYh
Lk+7UrfLq6Y8uySkgMpZzW4TOK8iNfJCWafRhWrHR8g1m2JcqTACzB3QrMv7GdP0
UpYZ32uwM8jGKE0P2jXd5Nts5fm4lkmU1u9tLT8YGL/xEWsC9XodGlAeiOXgIh3W
wmsjak6CVvCG+MPzsppDWXOEnaQQJXnLHgkUgrDKsT8BqmYivTqL0Ifpluo7W9Y5
vrVr4VmMZX0zRUUX5URwrj7jB08C5+yFlUYsKRlxC3pnjLdp0oC2yRrf3Ax0X655
xqo+s6KnW6MyTxZ9VZzsLjWxb1ZdiYWexZlSVmb+zXZV8mlvhPhTtuue8dD5J/6B
SX2LrX3D87n7PZ7XSZp4xXzXguo7f0Jt1T7jh3QA/aBn8Wke/nfuDp0A2uufFwcW
WnDnE229zG9I1PVIh46LLW0XkkJVHYGaaPWv6+qCZMiUTgcT1AaxXMrdS7OzhnZc
JGZybrHMAXn81aOGAEv/O2HdyRQ3fBtGDVOdxwkfFDRQ1vUVuY7VoxBc1d0dRq59
g7Dd8U7gAUR4c8qe0QhJvS6QXDgsoJHpFaJ70yt6P3EGuhutcaWZCOQevcQzU+EL
Vkwz8L4MhmTTT+cJ7SMs/4tJfvDBTiAqfQLnGBDeDj2Rsbp59V2f6zXnckf3g/70
JdKA1KTTvjq2Ml1COBBPbkwTNpZXQimt0WvGBPBcKrLP7cK6iK29LNgUQk2YRKXV
1dP/+7P83JTDPire7lUnZJM5K8stFDCQI1vPiQkKNxfLB39Z1uC+fxiIzXVvUkmg
ZhfEhVpiNR6UlrW9gaVf/0PZdrTMrN7Ke0BonkqxHxv5l/6UvcBXXOXTAJFTystY
bQkrRe7ePQxZ0YL9yDdPMp9zjgeyT13VxoP/JD6PkRayjUbpMJJaXrLYjdhrG4gy
86sntF1hc0qEUlJ2/YuStwCT35H8ZQ5SnmAo0EMyP0tNYoHVFr9fYL9IRJaSRw0G
1Mfr7LI3TYvfk9lLm884MP8iBVOUaD5cw7QjZ016Bt3ys7/mXuTzCe5C7uC8KtBt
AclFvCi3mlbPevj4B+6+nZ3+5aLV2BHVqxv1fF81yPUqs1s+5U6VUhTcva/NhQ83
a9WhsammE1lqhoH/MgJDQV1jIdYa/rPKmY+QtkiChWKIUxUgKGhZpjHPUx6r+uW8
HnXSF3nAxQUsuQ9RJuczuYkx2IgXxTOFum189MsxOXQCS+G3fbkmkgTlgD+k8BJc
p5kVfIk+Ie7xzFIyEhst827qM9BI/Y5Km0OG1U7/gSVVNAlnEyTRVuavN2AXl0gF
mdAQdS5YZi95vTq34RTwwifhwsE6B8vfNjZto2nToqJtiMrrX5ZhITWsl5DnPHnK
H23XxxxvE5JHJOP7Fcza4N56xvCpKgyi0GJVNbJfD9QxUgYxWlO3rH2E28YM+6g6
miDz0TvxVuNK7D4uQSFNFCc9KSk6KVG3zjeGHPS8NS+tvZdiuDgMsKdIdGJahtVU
DRgtYAuHTriciI3GiPedeIBOWyFl6YEm++HBFNgqQReAy9Ku6OGZDZLOVSNJV/YO
q3H6UyHUpAD/SO8ANHs2aYSNasSMTQ5WIQ1tpVIzBV6F5HycsmUFoiog3Hl26VL+
DsPJ0wGVPdojKmpHOlquiVb9A2nTQPzh7cb1qwRPpuwsCNW9bQTRuonV8w1bIyHU
ZwI8t88Oe+djOCeoGTY56mwc5Wy6NFziQdCBQj6q6wTJNPlIhExszeiANcZpuJ9r
Ks2seHrAcyq5Y2O8VIKVjuQhZh9ZJBaP3k1BEfGl2BymJop0SkIGRIk9BtRB5yIz
Ld+/WuXxHQAzIwxEpbpQ8MzhzYMIs6qpmsbhU+u9Qjo1wvVtmuTMDB4R4vU1/IWQ
b+Nbq7OkliMcElBmpTNZ4r1EDy/q1b0OZaISadsnOcwusBP20yu0YzKE+BnFdxCC
MFOWUX4D9uGVrxEiZ5VJ5Nw+evGdlBPEeiXWvqF47byHiu+GCVL8yc2o6lVFh1Ia
K4kjG0pJnOwDSu+kTvTkCXvWWNx6uQzxyUWqCsXoT6R48CzzUfkmglYJMvl2C7TI
kUN8qDyjxYbYy4OQkRumEVCEKBOj7VcQG1NWYKnbY+bxPzfF+J8QJGQJWDe6ESeP
2ohAHs7lhOmv3BG3bp/nmepycF4JbhA9AsTVNfDQ8l8cfpfvXdSq5fz3ygF7aVvc
T6jlYVh8anMPeTvgF8ho3Mw014FDncB/15cZZtpeSXKP7ZuX7Ua67QlaL4AfkOZC
mLOAWV5qTRdzuyrgOKeeuM8JC6QRrIOh5nYZq7GuU5ajLQvflOyiBewgTs7MVeSc
p/Az+DDPKfTk/7w2O0AF5lmn3rQhGxLsq8cxmb+PKUDs5yY3CuZfSGWRpdbRiEGU
N2m3GLWl2wHp8ziIRqLOQyGmcMOj9rYcs6THRf41+fABNLpM0AyzImseB4fYvuub
IRtnH1tbdgl1a/8CiJcPQmn90ARyyhKL/44IEAq8pEq9lxagPq66wYwW5H5dD0y7
BLQ6TTxjlFRvvx7C6kKeuXD8aFWNz+qTx9Xs780i4wj+c2vUQDfxW930P/mCm5m0
0UiVzBSZym80mxVnz/f7TIo4BKrditFRM0XZ76v+SPhLdT/0ich+kEYpHht29Xf9
yCCxGGGL8EPshx/dsqLor6GAxoHeWugYaJ+WRemC7NLWdEJNVuccbNvZvys2Lili
QjxYLTlYGgkj4rserv5FflTmPIbrTXL/HbFynx85OgQzR7gOddMi98NCmcYyjVBp
E2M/JgtVr8lly8aKY/M7pAT/zXaT4GWGiTPRkKX4b/64jzCimljB0PjkNezGAKXT
SD/BGTRgFaVUw3A41FQM4Fblipm/vMHScWQNxnM/VLNpTqGZMW38v4Cycp11CFXo
Ev8NvMV9RBvF5RvESCS/4IJ9tgmgL8rdKB3DyEFRxEPWn/cHfjbVOlM16C+1cEy1
fnMh7EXeKgDHXWVjTrjVdY+ZrJtx8wv4DmwmcTO2WDrnIvcevkBjDwSzd8WJ97G3
KmspQp0hIrEqPA79WKuFu0deT239dmN3rmvVTMswwQ6H3nfD9/TiY+lIqPyKRG8Y
9rZ6UWAtRVk4/GoUlNcrUedkI2xzZc9BsYT/gJk/6jLIk2eIuMdgK/Q4TpjJozze
0Hv2wOIU5xvpza9+7wXqX9vwC4oZjpUYq3WuwfB3CM32Jv+ssnA39rqsZTGQzsJa
gRFd70Xq0g2HOu1tuKyPZ0nXbyWHpbBsQhP4sKU2HcX1EhQxLY3Aa6TXD9a1jTZl
ZjTHywKXjRDW6hW+vUAXNoXZ05FqQNWbWgkWLBRSL/10zkkYsU7Rl4RoBJMJXxLZ
KxDRzLQC+bNjNnLrXsHQp2bhqSiWB7sTkzhH99qv2ST/LZjiqqMMqS5agkFbuFsi
AN1E+bMQU6wAn0ZVnwbncuBwsHAC9L1jmYer2XbcZOZ9SMiVmjkj5T2l/i3ZeFhy
IRs5GMySmmaUeUQpmXF3x+fQQY9VLvcMrwtgOC93tg2wNrDpp9dsCKDbyC4l43S1
1OITerIrtbzLto96q5GgUYTD8nqXOpnjSff9HMGvFNksdkylsde07DBI8686T9mp
h20LM3JAJLMbe2eL+zz4JD+cvzTVQC+oD8JgHrxS9O3tF+LsNLDWro2YxjKbWZhf
y2kYEAcNtIzllReQKpR1yBcJPQ3xg9MFxjbr6Ia47nWAFzuEvMy41+df4wHRO9tL
14hddar2AEuMZxSYq3QuR4NUgI/DOOxLIhh8MpXir3aHiJVnBGIxYtkIub1F9B7g
g8skeVyNk35tya2GecPwOaafvE5JvPDIjA7NeOiSq2l3cRTaM6slx0n5x0avo480
9lvqW09xU9ICizGxAwPPbPononERvZr3Fu0gXNX0WaF5qZ+8Hk67Vb8tJy3wA0/f
dHlHzw88jje7i0musVyKw1TCbTRcVbq/ROkOK5RUOpSi11HXrQ1a0XELsQ/6NYLK
Zatf2gt3EwokY0SLsJg+spsZejyngIiBxqvix18GGLI6PpZMKn/f56m07XcvP5xN
JA/AG7UnVIIMRqttQDFzdbjTatZ2QCpFvO2m9NrsL58duJJIzXiwmR0NaUEC9SPj
JXVhr0sontx81KbMeSVT5wHg6SIxK58ibiL7PRKk3thENMfDKc/GBxj1bsox+Wkc
isSM5v799UUTP31se+2d11Fs5kBlqJxQ1+OJi2jnwMbepigtnip73dtYFoqYVUzV
sKsze3uihzaGQSoInZbvjMm0LuEXgCyNxgtTjPF6/J6h49LNcktFP/47rGr18UmC
WqWCl4Ah7Z5QqRApbs0OdObAVm5r0Wmlf8a8IWTEIjWGE4sCDU5FNLucmnSdXvZa
CHfbPnItVRU0BpzxF9uDAR66JHNtq4/THGayh/Us4PMcodX3OY1kMbnlfwSRzi7m
gnKBj9bCGHiEmyjw4i3RNsQ60JyDpP+Re1atRVja55BXCuO3HO+8Oyva+QG5lSVu
y3HRBAv6Rg31Q8zU2N287mB0EHFRJXf7JB6X2fGZdg3/FIkKbPvdSJWTsmIbM0hy
fx8pu6hWI81Q8LP1A7blleVs2dn39byYGPJVMYHF2GkkEi/orVgbvvtcwGWL580m
bW0UQjL8vAmFGeq79jxlR9HM41dG4DzzV54pL4RXucPAG3fYNKrhVOaQlhQEyTqz
JZGXgr2qE+Kwk6G1+KonC+D688hQLGWuE9xWKeiKvOo1b5OhGH2arbn3QzBD4/TU
741UoiAHFbewUO5ammzRP4SEKkIFoZImEc2zjTEl44I19RllYmGWT6iThuiF03aJ
YvCwbz07pT9KqyRPcveiPHJZCmC+VSU1UkKYn6x49EHzE9CJH2l6bDkS4eXPHaZZ
4PWidyTgGPzY8iET9u4iY3NuKAaWPGunc1V1KWvmMZ0/V4EpaVwBqolQdtvGFUPR
/SXk3uGzTJz8t/p8xKlg/s+UlUYTHP1MvhWVfqRlrKaWnr7tvOZP7HZXGo8yeVtP
OxCU3PuawY7Kyd2c22/ed+HlnB5xVX78WIFug+YvZ9wh5I3ByRsG5a73Pvz7wIVI
/QZLGBZK6eFkBd4EOq/ROBIkA754KhySgx+T+X46k20GLxmBlmCcmvz9rAMEu5Y3
AyETNwnJAj+mxxg/gr9eAIPOlOrw/J5WZknrraTDKrRxCss1j2uOhGjnLuNVDpbk
oHcXP9r4DBxF9wxMbPfgn+DpQvmTUUqc0pOkG8WwjCehbXO6bvUOJKNacKSnhrxY
EWceMnXWJA6msXKMMlK86e1FmwafU84b7jx2Y2CH935IuMN5rg2FSwvlI0m1Qded
HT0MLJS4VmXcVsgUzOvNKhyd3aNha4LlsgzK6OZm1zvc3rdMQjDi8gJLQZf3mugA
d9kQyVODWDLPb3CtA0mN1MB7dopGgQMRewqxzQZlvL5B0/3YBcZvUgC3ocYzDvEE
Mi/U2cfJCkhcPaTjHEvZ1xMZAxMxF181FUiL9Y3bhZfdYepsN5eOARXXowvt4I6L
TN/SZygcVHj4gck0jGr2zH0rgYIMIFeg+fHFp/nVroIciJJ9JtWjzD0CfsN3hEkF
Mg1N+bYQHlxTxHkBm/eqN89BoeINsHItBe9SjI7rzibP9VL1sSQLlfPoGTCzZ01t
5tGUwY61ACPD/sGJfnf6s4B1FtuRj0qYoLnrtoCsq2cv+CoKz6x8tVDxoHsLUf5Q
byua6Zc2dZsQXLJ3nZe9pXp5SUTQUF4oESyw1s7hLKjdzaDyn19AwAmry3WhW0+I
No5PgUYUewymZKuy4RWLPOE/9M59RlXu5EV7XyWMTJnv49tGddbNNX0OXebh7GH9
ylyEQQ4etT6GS69j8czIruMW2W+e9ogF/7yZ1S4U4mZcNu8wOzN/Bm0I61c8PggA
zMAqDBrce/xYWpfN3yUtzPWeZnkCF1ECeEk+OUCIOCB4DL8vAhF7wrId3JzzSb/8
jxqe5LvoYp0UDHYjvVCJ1b7WaHWGivYBp9Iqwa3IPBI6rLhhUy3j3eh2l+UKJZUy
5njAOd8IIqucw2yVn7bzVEfM432PEKbcEiq8DxuYLNVWPcOWYMnKFVqrRbs0MfM1
2iopYmyR0NWvOWob9+abx0nBIIS8NZWjERDIUbIBo8MZcyRtOufdAdC7gdwcanmW
9YMUZyE2M1gsuwnSslc4Y8KKG1mz36jF92bWrAknrMtJaCNYqK+mjCn3lqLrwLjZ
Om9C1GXd0uN2Mw58BIcJcL5Z17dd9PE9czGa2Moe3b8eHf0ShnJiRfzYQ0RV5O1/
K4y47KxYNgqK+KVG9xt/wGe1Cf4D9a2y+0uWwISo0IkLE+4+mAU7Wzo3VN2el290
tQRR1NP/O5jZuPS9Wrx2WaxUfVNr2a6NxuMAYHoTaL4X3LkKHlriK5aUXmAL2kN2
+kKoes8B0GOSnPfjga6amtBk7YXi/mPRe27I3EQvEMkL2KIDc6cZDsUxx054Fawt
qiHWvp0WZONl0rY0ezMwGvWX78TW1ucUEX3WhEaHVFClRHnn9EO2kEcLeRXZ6UZc
k7T71PjphULunJPKMFIJ0OzlQRJ66mCRp8jKJyRXqtsMXw/VfpmsT7z1hfObJyzJ
V3fLNQ1z0zgs2Q+T4IgsEGoSRD987/V9/y3AleyQvM91tvf6rzBVjtQZN8NRI1eh
Y1pDlUgNkkevqnc/kCVBumAmOAgQMTwJl4EqyXgA2nrCAh0+09r2a+LgLXV0yqjp
FqGTn6oxGf+0pgw55i4hMpKJ8plCw3zK70zHS4ePeoXT4AEp/RA5HsCWK5KKoijl
msB99A3SL6Y53ADeEMWOtxqSExP9ZkLWLic9FAIOrNBJ8MgkPXczyyuFUlNHQQEX
BYB6FbCwZU2XaoQm9XMI2bBuVnoHjhjSIokQAPH2ZdWzzha+38RqBDUj/enN6gCU
bWOegcSm+Q9NpDwRXrgC9MsoA8CVELm9/ELHuO3AvRZnOLIrZkb4HUU56l01PtwZ
rp9Yw3W2H3BVJUHIZKrWKBLSdBsMB89KNk4klZp/Q0YIeOYQA+Pa6Hfw0A1bBDzK
yfIuApwFgqhiuQRStB0EXdXP6TX8xU1LCFD8LqjDQqtEWDx3+C4qvTJbjkBQI+NQ
LVY4qx/xYiWJh2qKRWgTUtGkZjiEkZSNgWnsihKtqXLaJUGd4ahsIun18Ji+UAZM
UQ8Zbjk5grPUvgGLxwhZsXuNNX6Crkt5T1qJXNPM7toKA4Y75cPKx/LXnDHSdVeJ
sCv119egooZBZ3y4WlWYbSjoz134ErynMqO4lthlw2C38BtWISl5UMOrEHY6rMP+
CLC7fFpc8wB48CrPdH9nWKHPMz2rih1mOhokv+7JUJfqToT6jzkUY1ufC8E7hl0f
gIc1yGbVPmKKJdfwPM2oAAh1bTxIMlTAiJ0pEx5WrjfMi7BhTFbHRYseeF0gkTBt
+/h3ZQ4FElZ25qhkiNycEMXa04YxcTrHOu+qOttHt90xrcKpNjOGeigYx3OsZGio
LJPU2U4vHepgiTTW1VsWhfaue5vd9p1ma69pbU7vWkiesZUZEMo2qVZHcgMhxF/B
hFQdBh7Z6mTWT8j4geC2FeZvTs6NlRZzkr5HJyv9O5ibhUZGoKiLkEY3LbogUDtL
B2WklRlrlCrck0Cg5maLysVhLcBjIDbynTDuzaD2Dq+9c4XRY6U4k5kfNu9Zgh9a
7YJlRGZZ7WPrwbaBWo1NMh9gHVxINy6iCwBd2s8M46lnQ94RQqTzuykLxi8wRkPv
D3FMGBRoCmI0li64IoUoqIm6bi++Qj9MYcb6IxfUEjqA1LFGKOgIV9v+gneHXEsD
t7XJdN2xVtaPGY0mrHolPDX9SCTPmvoCcxsIfmn2tV5PxhhrDMzX/4KS6yzEpUwf
lW0gvG+y+BdRTjBrk+CXp6HCQsgNGGGzCxzqs8Uvd+hayC1mlyUsUmeX++pOrnNU
Hr2zDWHNSdls0HQ7M5xn+IR0nHSnOTnor/uwBrR250aTIObrPGWOaH5cCGqSWlHZ
w701PDAEEJZBes63ryV2tBlzPy3gi6Y1/Gpo7XCc3ztkxzjUwX/jwLpRe7pYekNZ
E1irfMYNg1MfClyiJqNQbPnO22/SMg0VLngi42TXMlHwmyvAF+VjEtSXTjk2JBbM
r6tsi846r2WzpgUaqcvHkMHKWmmPRU/oSGPYVwUvGXY/33tZSMkJz5ooyyRXha2E
xC3+uJXhBHwd74ZO4r3ggj6sOfMVOIXRqPQqi0kX0+lnJBubIGKri68KTCMj0D32
7jCvSQZPRNEIHseItySB9WTlXBUyGUcvG1yUEYoWZY8+3N58GbJyXdeUIqKlWTM9
sjQRcgRs0HPfflWw0ECLy5AP/H2zazI37Lfr+oMm4e7bk78TpUzLqbMp1vjddK8l
qgjuatICfoQ9hvNm83MbUbN2s+EbRk4xWykmXydvK5SI/8WTGmEkT4p546zFVZUE
IMRolnJCNEbVCchxYqhKj1r/yQxibxwNAj2qY+aK2qqnMShTJ7ycAGagJ3UeMrjP
geOybxwHePmM8vozVeVm7KyIar7v5ChjTH/dKOWFjpyaZewwXkdCC5MPtCKNVwUw
60vb6tm/RsRvL6KknJgD94iieKF69qPSg6iS+A7lB8ylaUkO9Zh7dJIqisGOOnql
/KuUs+U3OXfqqR+v22TSZ/DBKBV1uEZlDan0Isd0II1hpzv3GFDPhyBOZd3v9HqT
8UAngouUfaaFFj40iq9NeRAMx1sMqA6/2xV7FIHqr0h5CLI3aG4cl94pwbYvw8ij
vTLLJfoAetACDtbdosslnptXnq5436Pde2NZV31GKtb3UnbdRoBTEKPHYfhRq6oI
cGR13HowGSCXhZsUqAfAwrOmWpYJAQTGyjsMdTH9BowN/bKPs4jxpb1/89Fe0T0J
B19nI+POljm4ts3BLwDmMbj7+HaYbxfvOnxZtTYwLMuT2TzdHYnBEGjrFeOMrjud
SEdMsz1VnySBuUrwhEC2Goou5FJRqOtqUyYtVhIj0S+UTReO/9Jkn6w1M4XBVgCH
qG/etEBXr1dpR/XWhavH1qm7zn3EyY65DSwAsiU0pZomElxBt4HbRZ1oRGUWZ5X9
3jZpbjCAv2gVR7GE7Mm/ecDkRqN72fwu7G9PpdeD8BkoyGC9dO77QL3OSkxMSasF
fvndpPrLyQClfYQCKCgVNe7cWQt0N48J97SItYouq+xO5x4ifCxvRWfBftgNV5bR
ZVG6oWNeM4GB2lzzXZpXE1iw+1dLVTLMh53jE/u9lyic0g9RSC04g0WiJk49X3cK
9c/Jr8gM/9E4WJdCgB8Ew5NH8W2hA+g24aVCBW8TiPJ+cn+r0z8mGPLe5PHQiCGm
7Fz+D7NoO3t4ZdNABq1uGTNrkEvxyiU5SxlFZpLsVmPqqbQGsIw99/y5hzrJDs4j
1FNlwsZQoLpDheYUvnsSclWVrwfDWZ+XW0lKOCa3uBr+MT4MGZea9lH+Y9Fi2JIL
6lqZ4+XKxENOUeoxfiSO09Xx9xklpYnSV+vmAwBCC5cFmYjGGoO+tpsC3nSbF3VG
YU7zaewyR31wgY9ZLp+9o66628AXGbkYjosd0APMe3nb0yLCj2GTeu0xeurKKiyB
J5HIIqP5fUPpl80tJ/9aTNZ7aS7VSgxhFCWEabebzI5IgR0sMegj/J3LSI26eASn
mlGU2RhFezP0bcK23oLhrDabtusrtl3A/EoLiazQJ2XwVeGf/+KQLZh23KdEuf07
7uRrCH4ot8Qsv4QylXiD3N0arnzujJPNVEXhH5XN1zZgkyCbOdVlZk+1e7ExyqTi
/VT3FqX10LTYxsc7FM14VHbUb/KeaCpnETXwpSC3jDSMB6v7YcpfL9EvFb0HeAVT
B1RfCIDFohm6AVjZVY8WpXMx+zEmfspNfPu6k1JpwiV9Ye2SjH2fS7csbe0XKJgq
5wOJq9sVnwoi/D6MSRusJCgZZOMxgnkmnSOtsfSHWfreXVPV7wKuxX7wY8OS094U
3NfkS89r9GIiPCsB7SZ3LwE4+rBumGUOK0RsNWBR+UinmH7G8qnjggvCiORxC/Zo
c859IYwkBabzS+IpES7CI1Vm3Dv/OMpdDvBezckFEWt9lio5V2b94q1eE36uOdhX
b40q9lj1aLhGscqMZVXdz+KPhMoRxjd2nqfOTNx1C34PMBM3SqYrMhlEypTEavyv
h2t/d+8MXdr8u4L/EtN47R8k0Azxl6p0QKuOQaX83x4GlYAAG5NXlIshoeQiFZxj
/gdIDzUzg4A+25v7Q8hdiSB7yXatFgyWXnAbfA1u5D4NkqQo/r5XAv/4BqZ5eUQB
eSqWVL5jTaMVdmQiZqj+vtfxeVDzZ1kL8gWM7oQrn90UMiS2Yq7ZO7iWj1Lwj8uk
epU/tskmvDihh62zpwtEkGDXVHshe/RUY5rhCvBarE2P+dyd1me6FFMN8d9L/i16
mJu2x2hdMDL8GWi5yoOX2oolHolF9A4A05EO89n412fYFxWHR4jqsk6hjX3HiEXg
5dSiCWu4tdvfA1/wNGVI+4gemRBCwSxSuITvswsjvGbAblMiSiMaP9P8uDtT9fbu
crhmk74lHlbCfvfpv7KpivETN0ZlFr7VTnKymUXtsD/Lnf5pSHtRlPL6zkYT8LUI
j7dOH6qgGHH6vL9d7Au0d0D5r0EI/4ys2OqX9mgdd9Y0ilfeBC34zYYNlsXm3d6a
sE8qKmKhEY/6GEmhR2V7KJQPN0qKuAsq0WCwQ44bEEum3BMbdkMKLBSbXGeiuoX0
Oq6Ypux5dvPMw9oeZ8XZl55cMe8iL5JXU/8mpkoWXwx/XSqJ6FQNkYnzoFTKW2BY
uAgJFFVuNBsu7eYT/tHQgV6nNxN9VfQi68Qb6fuiODc3GXB7UutDoSKc9Tbzzvi3
FIhNETUWXg9C4SoQuQbLYcAMpYdNjaBhT0SUVoJhhPJjYPecGxI+d9BeBWqVgSxw
L2S41OVNGZrI0xIpoSh8hKljQfYltd0okUK/iPq2V9gLV4JI0IjPJXuwq7WCcvxG
bXgIOcrQ1yHLskjfGxKhUZ9Gf0oF1ZRgvMs+A/37k9shaRbZH6LswdMh2sOfA3p5
zKPWswkIHDnMqHOOUatJQCBDhPG6Tkhm4zsvteaVWSAWlGzjCSbCzni2zqjybhVM
9nD/i3NneXoN8KXlxlFCZ2k3GUGgD/iJs36S8RKFyRITDDB0UOMkxQDwB9Xd28JQ
jFtM8nr8AKoE/BXBpZLdhl1aKvG7zbiLybDcHBJtAIKPkhT0ST2FVEmOrJgyq5bw
dTbUapQKXGh4fVJUDMpLFnYtFZN2A6VL3qdkzamJ4V2kPxtxl6GcTetQ6V53a8L2
a8dHH5vOqRwSSStS8NcJdRLdYjHpmiwpv/4/GwLgHywhTZvnDyXDcNJN4i+JNo//
ZiOGFYm9W5zaHJQF26NqYD4Z5d/867AaNOnTyO59EImyZEe8Aacyq6A/l+RxgwPZ
JalIi7y21r6/kqLFgnH9VBBMMEuwGrQj15b1jAvE+szfd2JvbqUKFW77UxTUcClI
ce9kx0am4kzrE9YDy0LoBc7pTjQpXKOzlSs/4mcSycI+cbkGFYnpiQUHIl4RhMw4
ARS8ghXFpZGxTEuscOKgsv2l1Fxxn34IHADHhi9RWxRxNl6h5+k+gmBTBhfKoZfa
5TMV1diIIAH0vrQGsK8J1uSNGT3+z8LQYg/eEaBlDlsu4Mu18c0Jiv2BfK08GXzg
hPOZMPKjr1ZsHz1D9KyWPaCPCMpujW+pG9yfeeVSFRMIE9os8SeKw6NZQ7uyRYoh
FpvO8D8qcC/euf6U1frN/IkowBV1XvoQ8nNuqX/RAyTfnOYtg6ItCSK6/iwFGlg5
VcUJXHhC2FBpiEbN8SkLTbdCTKcZ4Xs1JCTy3S8myk0th8JsrUrKFqe0sO5UiM+Q
poX1blclG+3Sq3zlfOmrXS3c5bqv/CBIpYgW+h1GZUPFzhAM89XZzkksxOv5zMKV
HxLfUihz1RJCEJyFHHij7YVErED4ABjMno0SK1PAGBpI84diMfM9b9sAC4XZ7sEJ
6CdfoPAyL3CjFZOiJ1EzVaPCrm9i2vP/lsWdt6Li5BMRf0mA8QkgzqTkzzd+mBXB
LeafEg6/TvG31FW2yaOTg/3mvJLeoZAbE5y9BB2w2Kyp/2iqo7Y0sbG2A1M6eGze
RIsO0VJqoLFO1i+pwCjFa+kpT5D61TeQE8h7SKWeKvxJFpPgupme/U9IqgP9Fjxt
bgTOvvnKCe1wJnbZ+iCQEey61B7mePZPrbe8vcQv+S1igpvm51wpWOdo7ejwgTfz
XrfZt3aRlafXBZiaeMfM2Q+JsuJ2s4PPefAX5EFbMnMlA6XYbEl+diWhr4/kTbV3
Bgf3iAhJudRc+Ku0i2QDrv5PejL+nQVX72aJf/V0YsUrKmYOaE1gxxjwyMXJaR/e
VDvx8todTMZCcqKbXE5u9xjuqsp7vabRpyxQiQRKshDc+2atfPDp9qc/4jVUFCkL
0KXFsURrg/KV9qJiYmxNReaMF0YNgF6yUeWZJINgz+GrVUiCZwoIsVMA6Vb7cvvn
yfuQkYDr79khT5bc0y8xAdXLnGz9VICsHATCQ394kV8wKwMoKeCf22ik3Mei186R
ZSuluaP3jShZFH7vSkzKHaeE5q7nDZqp698u2XY/Hmy7p3Ct4dgAx4av55DTnMiM
u6BWTzKrJJiA9uV0mNlXQduw4EPE6W1W14xsLUHtjPq00HjQKJrK0Fxew5nIPMG1
PDvYHj8i8k54uyLQ/GU/YpZZjkckucoxoNZrZVjHWN89XtP2IN4WvDiom0AZJQ5t
qfunGhg9uamFw6yUcpAnrK0YMQxlJ2uz81ws8SVWHQ70/K35MTW1+OxiLlfqycDR
tYjs4s53TGFswWGrMtEy49RL8Z5UXg06YcB/Dk69Cqw+459YnOxtWRaACY9itOVo
4DNgqsnvd3R2cTRwWJOY8a+3xF6DC+i9k8Inc7s/hhq3u21gbB6SY+o7MqgDfBtx
KUp2h+EW8Dh2kxdltLToi4qIyu9WPlH+Z3LOvjIEMAxpkDOpW2RE7pl+UUHzRdYf
O8qMhio95bnaPWJ5QpefxIKVxU6kY7hWrgPkgs2clmpztHjZuprnKD3BeQ+jBpEd
/So8Err6Ey3GY7PjGauUQCzTbwD7uoRlPGawBvqHvMIpkJSoddi7/rz+4lx6jqse
UrOlqBRLwiwlNePBcdJrracz5jdQJWWUsUVXyf94r/FSesFQywJtq+pcv4sgz1Jb
sExAfZOVlo16WG3EQO1WB8XyKyMhoqUd2bhOwpWcEsSoFcj3ckdLRIRO8XSbuVOi
n9IeX2spnlQyJ2v6M4YYzRECwMCjHnwTtupzTh08p1OxIwg79AFrDJso1GzRrgQI
Ym82mdu5+H8+f3tgm4xBsKyn/qIGojmg2yPVuZWvjRoW0upSFxXcIOTmv97oaII0
171GAFBO3aVzOehyC8j2uYzUk5n06YSPIq9VisSyDcotSQbHYBkyp5uv8IXC8R10
YDdiNM5kq6Prl4AaJjXQD2yFP3BwrxEpdT/tU2+oxBAm4oFyfOrBxko1X6TiwIJx
QmZdognwzwdngXbemdV0BcR/ejbkkMvrzEJI9dA3tFm5eQ4PxaPAdZhUZbHgcZd2
Li16zuBgC5wZ2YGel/Pa2r4ZHKng8x8Q/iSyFPL3ZfEZib69cv+y3fHKZP+Bcn0s
+kRS7wLPBnhSw7/nnIv0Gp5MUroKTxxsvUBFG1uOKssNkd6JgQtSzKbkJy+D34uo
6WV+EjUS/rcil5WQRivd4rfx8z4PI1NfdDCf1JCdROM6QqRk2I3LVayEKANFj8x6
SJCYrhsm9hDZbIsKJ7m4I4IHJxkJD+jMZ0yyeIxXobHyNs0V2wRoEeOflGzMX7i5
+4dn8mVjIFeL+DG0NHi2/v9HRWBsw4EwBJhXVwrxj/drJe1vgamAd358VX9UC1PX
QMy8uMpZ0u77fL+ySwQujhKPTDT7weT8dRog8gIpvySycJn2F4T7EKRN+7AKJpIh
IgO5Us9W/SO5Z8CgJrKocYQIh3SKax6geI3QJSyeVm/GCXBWNW+BuqIUlhLFgU05
AMPC0JyFEXMSVxtoXPXPcUH/weIVe0O1mhpObQNwlhtIwM3QmFdTBn9kXEQZ3gvH
x7364xsrHOBppFCTcHcCqwplJO9vhOMEci1lTOGxaXaembn+g3y86t0Y+gUKHN+7
wfbxXzT35Fl15kGWluz6pRUJDPOXUsqlKV7cCR8iCum54c0RRrN386rr7PlJ3ldS
znqRAggCOKns0QXio0rPEn5OGJvsOMIyuUWrKXOG/8a6m71+sPc3fRPTbJE+xAbx
Yp6STuI9yLxOYUCQ9n3pCYEG5RzgwR5feMZhknyvPK4JpPWiH+7cqwVIkEBaOJJN
aJXOdQdt/2pFoBQFHxXY30bxbqlcDjzI1AuBFrhXP68B1uj8X+aTPZ0GEaUr1t5E
AgBZG1oEweMFVJqCGa9fKJiCgbMx7IsJeiC4l++hH/L/+J2v8ZeJNgr9Txm3ey63
5qGr/cyBL7cgeTfwuTKVJlq34fKLOBjYK7pKpTc9fBwSjNXGaSV29YAw4OvywSTp
pxV/SSdkoo/UPGi7Av2CsJvI/y+3NQOC18/xjt+Ea7hieoa02uaHRlDOMoCOYoLe
glTO0Ab9HGdm/ywcndXFOMKNdXXq38H3Ls1z3061blYHXZbXlKzU7FYPomEc7b+g
dmyFO2pPgouC1Vnce7tTH6KUJSXbth8bDY3QAdHE9xVOCSlLPe6ZtooMoZvOmtHb
A8O6Lar7PAsvobgHvNba1KH0TgwtVZT+uK/YsCg5a/r9HENOKm13M6TdNsh/38kd
MWPBfJosarHFEFQoTik18qSoe2YYJY3vE6gZNxK9tZfDrZz8JL3xyUUgVGtZmMAM
WHk5fqVthW2ZlEHp59FY9WPa9rngc8TY54Jp8jLM5wvtLEiVi5NX1OEO2ohoEUK1
SU/cCUxtnVfyY9qdaKasSYlF4sdTWKMoZQRF7nGIbZQDVCYpTT2OAmfxXoIq2EXF
rrKiETdFaOupgw/Ug3ephek8E/wMliuSRdR6/hjyKYtt3ue5wwceyCKvfKVgxB+Y
BRC/wS5q5fwcfoO/vQhkwjt7e/IqlBJc4JejHx6u0logTW6G9o4heIUmK7GoXbGU
g/YypQVVbG0omJjZZFVxR/vyDs259gHSXpGL/vUy/0Z/m+xw0FDZ4DB33Ot/wTJt
JEptRQAd8TzoCLbnwGVoOuOoJIdwkwsw3fKBVoJoAsacKqe6qwgMJ1hPXOqkVuWQ
Yj5WPsN/regY85GwR1ev1n+SfGpcdJxNZUOEgYvSShFDoGoPDteWgiMhwqb2ThzL
st8bGmGqM0F/V5uO/++Xa33wJXIpDivZfjbPIjud/zgGvdNnk5NuOVl4M3X6oOgd
BxaDjWsI1V2cGG1GezoFmgmbQMWiA8F8TdPNNWMuv2a4PGSGLhJmROCJS3d1/6+W
bXX7t3CZFm2SJkQJClPEonCTmPslgxXcR2l0GF4iHnZDQU+lBSMlzXKNGcvBI/CM
NP+1cMAWjsaZzOugenf6Q+Np6EAbKd1C7sYiu9JwEyBbpmT4G7I3Arh+ABPanSxu
bqkA+7LP0Rq1OOIJGBWdU/jApBd/lmY2+BrCrUUCxcmileKMNMdiFqvqJm1hYFPO
0q2IDaBuz4ZKdAl6tHn4JBui0hRD4kwkSBQjsAjSMG6c9dkH0U3DkPQHzu0vedOt
NKVY73RmI5CYzzfF/nIZcxdSJcL4XvpxfssnOhfVYpRIZIQKvhf1RUIW54bAySCX
dmzCDZOJhUaurZZZbcYX2DKsYh5pfWWCpqtvQzgFkokEnbzhCEpjr/zJ2VRlqKNv
KqcJeiGt6xEiDc1tHOuOCOdh8byCeg3y8zbyHu7fPQXADpqcGQWeRLAd1YzcJE0d
95/87TLz5CXqb0EXKN4/3cE2i7SBS4eGRKrPp3Vzf3GRFe0Ai0R/4aH6HTu0lYqa
cyr3edQfEOpcQWDy4wgfBPNLZ8sq6csVU+K1JWFDHUYpyEmaiHuW+i7Hl7ZJCCOn
PCxbgWWaa3dfJ2164Y1tOY7QUsmZZpl1pxbiBuHV3M1h4i2TUgbpxnLCD1jkGAJS
wy2yk3/bW0boZZEGP2g+wDajP5OYwdOQzzVOXj6mLqhNnZovx4i6aWN49a+mhW2H
RJiZng7+zcQ5vZWdwfGEBtIXqtcYs8NRQNz6kEHDLW8NqQI6z8lO9pO9PRlWe0Zo
Vh8ewLHmRoRFk9PptWa5V+PaFw4wBlnycfkjWMmw1WgYgaM4jR3p4sE7Cc/uU6LN
aGgn0YWIk2SNSWPKpm38nEYNovZyWMc8S6bJWdqK/dZeXxduRdYyEx1c4vFpyquT
MV9IHtRVUCw726PqWqKOCMemT2GeJzAlEF4KtFG+fpBpgWEO8mIMWMnk2eHOHDxA
XhbsgGNk46aaFyBxF+sQ8divp0AWjTCNmsEVlDEcrHyArqAimwp7ojHJ0Ed7qjtr
xpe+qDtIosIh8EdeiS0VMxZgS2IXc50hVAt3ibBnCb/8UbgRsA+5vsNJ9oEJHK8F
9Hds913PLvoM+BeuYVduCTdaKUZp02vU/97vSrRh5Ktgg0V6H4NSnlpio1INE5LS
259wcpCin5DdnBy3iVO3kk7AQEKjiYYI0qGh0o/bGeyYBUJXlyXf1zJL47gZro3D
T3XGOmqy5kAlWpPiltMqTtdXgONjr1FG9+1CmKSvZLzSZNBdNgABdIKDhprQ5xD9
XKFfJHoZadETo9CbrseSp8CAArMAbNDezxHcBqU9zeMbQki6hgBMUaQlVlDnQ2c9
N8f/I9CBDygCA7u+L8GhUosOBVMTWgNQrqmrdgqJMVifEq+j3B10QH0J3SdfgkrH
N+J+vJ+g8sJYc5U30zUIqPfjiiPZRvAb4+5ONQ0wwATZbKgNSQ4PRImxnhsUJq8f
0V4XkYMjYZXTgX04U77sUDoSrzz3hhUAGlthGPzQuxI5xpR9Bd5LhwVy0Lex+/XU
5SCSMd7mP4LkKVHKuQxyzpY8+Fq9RTR7PIMlQcGfv6QK/gXdKm280acwLzo0jUn9
qa9OoH3naichB+AVpJ1HHiHUn43CLAhL+Bc20eV1Cpc+swpXTbDEaS8ZyZFKXyW+
9SqaQYaBFtAnKO1sCN4hnvplBGFGZgLywswv5DWfPKsSbLSI08z0oJaGcgXouW2g
fKeOo+rWkt70o1l40Ck5ahPWtnCSitk34L61i122vRdr61x6DSL4/7fgaNLn/xOX
8kGCKlTHRtM/BUBNP0jQirORcSf+O9l854mm3g8f784lWN2blIuOjuvvkgeu7Te2
6xaeJcuvhptEANHHgYR5MzsbD2fGfMd9kEqzov4aefgkBfQe1SS7dXCly914cgI0
uCgY0w2vEUm3y1DHKNUjFUm6BA2LTTZAlKgAUF4lN1oITJKD8owrG6ukYv8p/uXR
bkqR+06hx80soubIDopY9YQKMHXCtUqw123Lf1euLrHuROeZ5/8MPd+VrUBQdnTW
sd/f3RpLXlk1wrg4jkPmeFRiXBnNNa1AeoOizCX+aV9lHMzNB7vSMsrVEHs/kazW
V3aVwKTLm7XqceIPqBpVIt84qVQmsCMRHbHz7pTF/W6m407DA1j2Rc+59/SywxHi
yeqcZLZvBYmDYa7/GbDT9UZ4neKR56KZHgBeQRGVmsa6W/pTn1O6lcfugctK7pir
Yv0p+6l+FSoihPAHQut0zJw1QGyojU4ELhJb2F4lJumBhZnb/kvnNnBWl3xikBu+
QpPry603wziOVaNXo+I3+h1IV6OMMfGQ2c6yhVkjWkIazZM8t2HD2mbpmI8JcHoa
gfTtNU3aY74MquA/EDkkc8IL/1NPtualElsj2RbWeMfQTUcvdf6GYRqY7+uJz5GM
3qKR+zemZ5qXpHDd/xwIGftoGieFJa5S2CDL4heid+tJym+xMW+0TrSVcNreWE77
ZurOjh4KBo+cf0G+Y2bZTmekludWkXe3ah7fB6YtGHu3Izmhpd0XNbJPZLRAB0do
rC1RMeHEMJH2RwpF4jvLFFLEVcq57K5qbXnMNe1VmppvzQwg6MnsABpWWmJUYBei
P7GWlU8DVx3MPsW1YFShxPGyyphtNC6N0PsM1TP+hr7WQRsZP1IfbLYGuEPAGKGR
tLoZu/nPd6g1u0/HprdQQPVxCy1txVyUHws9hIIqXc627X+TcdGKPAuRqfcLmTzE
NlhEfiJyBpaiezZTaPF1EnQNnD5AkfxoenX088BL73avRcJ68m8UTJSL7nxbIhbR
7IQ5vr88RnDU20FMEk6EsaoLNW6r1wfekVgnUc/5M6YF54OGRJ0JDP2wX+1jjPHc
fbxxpVmJ8o6fQaemBE3oGjUO5lvIwVj+a1xa1j23p38DdpodsElqV8b+o4R6vqOg
20AQKhQ7KAms+ERdR5OFLDl2Mahch7piaeP+rk+IC4Y3Tx29lFdpGtdyUpggH9WE
XD4jXn60lySxdv7tuJqc8PBvwnCfWGJOm8WUIFGeCLU/o0Z3kn9FTMIY6IoaQbAS
ErjueE3pFr6I+MdebHHCdvw+ziiqABM+kvh6PmKWRvC+gV/haeDsn2w18LotE0PM
Mf1+rpJb0vSOrDXltcMaM/iMixIKkjYs1JN5iwUqOww4Ch1wgfVBNwx0ZdkcPQpH
XIza0Z/FNlJZbOmjsGX7GUY/1czdl4/o710BBsOVfLh0YzKZ3/ET+9KCZ9uQaljG
GK4UL0YopstktcPvnc6U0YSu/NcSz8Oxyw9ikWLp7wd254jZqCoBkfY8Um7mQPnt
5mxivNfjfDTFxUaJzIQbesi5QDWKZky4z14S6nO800vuvdRnMm9wTbdFWWss7qhR
ox1gvLniXYvXv254vHc87CurBs7EUgkDNFHHoQxfmHJ00PI9GphgVmxK3TIu7wHV
+wqNPAV3r4nsi2mv4fSFgK56VtA3sz0DVlB6rFreUctfhUz/SpUD0QYdi5NTIvpS
WkBi6BQijwKT8l+3jcpZG9bzfC4Kg0cfgdxCmBPjEMVdNPkPmb3QCxRSuNFAXZJ9
P0IGTVduXFi5uXf8qRumbxawmYymDs7uin75+1d/etXMSwMPV2CrkVZzaRCL14AK
HZiZz6cvHmAqiHA4nE0zwgQlFArckOT/NrSlliwhTadcLecVD9LeKjj/HWm1zCKQ
4pqBlhm/bK52X1nO3BgACx0T8He+v8hebiJqAMXavSuThux7dEQJxlREafPWh31R
iyUvNmObGgsojDwTXFNh9M/x6q39JA6fI87LH6FA0lkGcf3nYdUxtGn/ksXwelg6
djZUNBBO4yuOZGWlkkEypctbpiPU4bEWztVFmPCdc+sOdMucPQ9Q97N9kEPTgb+8
r/f3HiT5pQ5RsLkHt5vwqqkD7rUrHmBrNrN1aGWY2dr4Ujiwa+hbnuiBqu+AtUby
A6CeHt2BxgR2FL0L8mAR81ob6a/kvRwJKZZoJ3px4xY9JY3LMvqvvKNZ2EVSWyhi
D0c6f/ZAgRt4bGhF3QwXxoixZKVm/gjth/XuwQQDuzLXVQU/30hL126F5W/rlvxi
jnOTsHAwXJKqY/EmLpcmB6mR0uTzxBZ0IxoURPiRROLFEy1gkNILM2xCYUTPp47h
jsvgLJ+QSxuS2ftoPlZcenTUm69/GSGAL0zq6Qq6AZ6Io8akFe8tbfs28N3BQySq
LAqutexs3zATviNLUvS0RweyM/luEABJsKVAYLolHc34fMQ6VZH5iEaHFxMhiP22
/i+x9X9F8RBvuZYhtH20apb2K/Lz7UBWuleeATYTGMdlj+6IAVMJc7UOznaAWlqF
RO1ewPk5Yo9gh/tr/SGfHt5YAnIMtIgWZJb6icgFGz7XWFwfiajEWjb3EKU9A8Oz
+NXHVcEgjfoeKM3t83g9b/aZC/VOAlTvEBzAyOjN+TUHNWQlQrnsiq62iuaIVcyv
XY0hOHlNUaUxQtxj95qZin4sL5yHxMyYb+X+AJJmrttknPn9Vc4pcyindKYupsxi
iEGvC4x2E4j9WhohzED6VA==
`pragma protect end_protected
