// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Re6bicS7heAbqQ+tIjqVDe+boZxs0FPyb3EbPENY69O9FWBWkeJl+VG5WF0KTEHe
5UBjCIbHqRfxVq3d4a0JNP5b3cFwU8CYz5QIgP57ewbN9BK60MmfWrPwR7SU1jta
YtAzkBgc+xuUyBrk8Z+L/FSVHlkwE4FGHEfQInihiVk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30288)
oYqOK1/u9xsTUIqjFXQxHkUDz0XLfkSn52f16YZGRN3R7lXN7MsbAIYaTrfFNu8f
IcPH/dzOfKurcH8LYChWvaHOyMYN5FldxjL/Yo4T9BCXwZMckOznp+HpepYzPMD3
zn6tvVm4byJbZ6vfoSrLRZAk49us6Bce+JGDzVWuHO9+F3FmrktQeuz4I06p31ZF
x6kRqdD5nnh4ofAa1PRDs6UOYmIYgmaO5lGrS+6ytRr/KTrTfHP3F8nAk4CF9gZq
8h4wwONj6Rtq/ht5zUcyxUHLn/1Q5MXY4tNUvd3Xqz84J2idq6rbsPj8lmy5N9+W
qgd+5bt5NQzjsV66ByceXT1IZnX/KpRBlORaklXGNyKXzkMkbV6UVuzor+7lwBN5
0MJKhffjJdswEGoX/boBUgHsUV5OuM6ol2IH1zILXreeVjJfxTTpP3W7cegq1rJu
NpRzL1v4xlsUP8mCG3er6oleefx+56JJS3cvO7+R67s5wnvu5giXuHCf7ePzw8TK
KILzUc0fouonrSgmBrKqv1lcfqwCgV+eM8WdwPo1rc9yfxRkdtldFpmEfQyk1flT
KGsdUG32DAZE1zVpr6ptW1AlYQ5m6hC5kaGYktyQndvxF8jBLJo91OofeYsrr6Y5
l8f0C7Vh7DblyXIqnIZszPF7kuKPWUBSuHE6u2oMYHutiyjAgnsNiyAlEpb06lOc
APxNeAUuXgmPCokAQX9HCqRGupZyBb5XWXoA0Qow2txRVeWE3NbdAQ3Hf4Uo4DB5
fA+/79fQEz/jttW5VQNHHgeQrMREebb+FB6ZHQHdtSzZdNMNH1is1Mxbu8zmiyWu
J2XQqZtYt1vK8N+rV3AykWvVAxbls8UcScPFq4hDYzGAx01UgrUOAeK8I7bXszUr
lekGZEcej0wsjzxO4D3Xvfa3bfTCdYoW+0dOXW20c+zLscsvVReaPztmXi6cMbnV
zwyxB2jhYT/cctzRBYerjh2eomry8Be1YE49NJQ/QiOc0sP1OqNQK7L26P8R2eT4
P4PDDoS8KDVcAlKWwmf8guDgi239nJOa0wjXBOLrrlbUzUKIbuodMF/QQgRgDbbP
rQUjxUoS22BH7FbH6ip8RTncVjkycwzTUuZsmwAYRuMcUg9DCEfWZOFVJTpELs63
12ZOHHzW/NcS8WVg4h9FBuSISkKN9aqpawRTFLvCmR+yh/PkhuEnjiCuOnxAqdnk
IRYM8tt0b0i4sFUun08qQW7XgDx54hBQqTk/iNLYVOpd9V5pYMwnDRCN11wV8Zde
IWnSKcurc6xRL8j8cfJp41/2bTlGWJV50ugXDXGeztUq5Ju59lz1P2FhRGFhT+m8
pBKNDtqfwdXfBVZmx/qkyKhgzYrTXx+p0AHmfEKWFz1baNL3H0kjETRYKLxl0CiM
lfkyUKIe3FvBvBfCDsRIoq52C3B6ir9z6TimSUNwNEccH9PmoRyTRhtZ1vtZpbxJ
Ttmy4YnJeQTAKypzBeBs9dxEhmMxg9BU9iRVl4N0Vyf+vk8JYSUIjGuIgZh69JB+
bhCSfl+Bm7PszUk/smppJgpEERQz5fEolhOEuQa+gt6GKyUcbol919Rj1Lj7gcFA
jOf1o819MvVwOCS/2jF10vZtUHdqMKLsK2We4TlT06RxvkEfcTiCxc75OtQLwlUq
CFxt+r08OJqU3HPXqnunXIhA8lXurxNAQZ+vEt0Vvzex2fge9qfhgprYXGZbK5LU
GYf3Z2M5eSd1BZtv1eqTS/p6El5gNbNqzDu0PX/uPXV2zRxJkFWaJmJ6EvI5UBLw
2iXSJjLk3VQkfv1/77Q83P+4sqP/GV2+yNx1asjvV6VwxQZkLT5yCqBKzbavKvap
5deunL9Y/mFvzbaBJcsoH6TXsiSTeJBeeV76jJeYvf9fW1HeTHRhsGZpD7f4GqEO
nEm9utk4kAnit26+LV22Kr5gLzIB0qTmhWoiaOSbi4xpdnctULEb07EvHiK6lM60
o0JvgTymme4ALQ69HAD40sQ7okxqZMjAhP9ieY9hM50BbQgbT87HwiCkl8rJwzrq
KpB1HX8u5I/EbIedr06P88nsSCqi6ghFiGOwTXkjPWHAYNZ2lJTlT4FWGsXNJO1z
FOxk3u+BUaiBVZItIhQE1zZHgPLWdcAdco5JyBRAnokeJn79rwKW0HS6iBjVbuFs
2w9K54Ij/hRuhk5CJwp/+cw1fONitN9CTX4flBPxUQkl3SPAINiAYihjsxllWnvV
g1BL+SfR0BitTHV6F2Idab/Oq1qcjKqXUft60wH2vv9Z1HGIQfSYK9VS6f7G3A3G
OOEwtzg9iVkCrDgTmn7ZcMlxNWcKgYrcClDB4JiMHC8gCsqXGmVCM1+Kw5Dm1ddX
YxCC22p2wk7g8nqc60xSPx4jwqWiMSS29oyj7TLpigCQ8CQxxdGekLqHMwphcvvv
Mz2MEEkg/GTehhgotkuYC325Y8fTN9+1IqBTQ+n5RTIlFcuUyaMiBHTOiUc0jz2Z
/LxN5x8FyVfO2UheMUsInX97oVIlP5HYTUiWcakPqtSe/+i7n3z/mNfBct6K8gyM
AVgIiMjvmdQ1DjR5DnhPpXy+25P8PdhInv0JOYdkQJ/FwVatKW0TvWwaMcpYB64J
kKhzPCK9qAx+juupZDx2yvpqj7SmNKSjnmx5tsQaqpCzhf7cpI9g1EwebUmntyqg
LQWyJImm0vSpG892XelJpwm3CRPqii2uGgNud7LtucCyQ9LS982YdtuMsnWUVvvF
WbI8ndPFwYNCMBN65po1zmGndhgskROEyf5d3WDlHgR9v1elzyP+1vUxzKf5G9Ja
c4BKBhzxgBwLBlwVLz0exKI/HVmxGygZLpaedaUMZHJ1mmwSyQC6R7xHHxXtrOoI
Qgx+3joKOkROF7E5sLuxnl5bvkTp+HKozf6kogfZTm+6XC7GXZ+WvbzzeCIFBkPk
5iRBrEO2iz1xrKtJHTB6o+ucAcL1KkshPyimrz8LuzhXH/I7LtFwD1wDGxMDFC1T
YItB70B0k3+ckoA42aFELIsW/Lyke76h0Ug7TvqE4rlO9Mq2ZA5961mtfZqFGIjH
fOuhboaObqZFym7GEchy/509Cu8yf15T2xzxVLqkliT7NpoipjgV9IybTgq3wKXl
JuRodnaGnXZRX6Ant0S/bCWhefiNBw3HZutci96jQTMaMCZmK6Ge/8n4NhNbozxb
v6O4ETgOE5DBQcXAo9SDoVYeTCLrHtKSYAfG9+cx166h5pTzGfumvcpVptDFJ4tM
QZDdjQ/FF7zb3RuUcU9pDfMueHe5A7D/AWVq8E0xJRdeQRrgwU59VrgnmcIt6s2Z
/E1Ni5xFC9QqWeMKaADc3/jtDhrTINW6BHq/XDOlkGMsTYRoXIAmFYik3pFB4hl6
GMQleUVmAqOAKKVD9y8Nq2oAJgqctDG/ZSGPgZIgyrQQ/0IzAM2ee2DdnC9KMANm
kBYhB66aEP0oC90VFhObtqD72+wFQSfSDvy6PTO53DzMYqXBkJAtw5/9uNViVUEP
8BxZeVB2A0uS5Xb8PIakTqHB+ODzM8U8EJTPeUhhRwYXqFTcbxWcpNPa0+ESBMuj
h/4uUrjhtiNW1IZNfemSzI2eo9MoNFdEz4Pfws3Sdp3Au76Xhk/Dm6dJtrekoFqk
3ampNCl3KAw0WavGjlN2UCkJPnB3qVW8Wli/ocUJ9dNwCEvqhfy8FtG2ZchC9mdP
Hia55MC6qi4pvzSO1ByJ/88mm/SmyWfNB3leolbBcTpyHsF+35dLOO6OKSjDr54S
rDUv5oO+Wi4t1qe/B+LciujWl29tRh1nUcKwM3zLPWov1gKOvvAlhXL2EQqHhO/U
o7iklHNWuGibqA9U+PLlez6oWd6O48msiGnBpiM4kZWgYEMr9scFfA36oeAvfKn0
GgJFI8YOMGtyE0P22XR0cDhg4BnhU80RGJBX4v/qWtqpopl15lZmBaBUv3iLhayS
f8FuZhAgWoj7UfGhfTuvCWF9dLFPzZImmIwQfQaeBLfxrsuAahR/gM71Pmf5+2LC
Q/TWI58WNegwPsCiyR7XSElBq9Jrs99xopEZ+tMBt3mL354GLDR4nzwFox0/xmm3
UT+IESWafY0K1tL0R8x+3RHgvVOSmPPm8FGGNuekDlnHz6g8mH63ljAPph3gVs7X
97syJpqh4CqMAX+5ndByrdoMmcfO8eKRhf4pTPRf3qpKZmQIvuhv4p7w7kyxNcu1
9+3EAPGiJwbfsZElsggqtm3Lk8LYp85elL59BzAaFqTvjAlegQs8RfEAa3er4QsA
9NvkGS+y5jxYeE8tdHNXTdOdCMxdSsRFR2ioKs/9KssmkeG4Gl0Zkn1XNXMGs+mW
hsL/KRBdQXvBpDctDA+1WKafl7DZok0H6xr0DuS1vCfnCAlmhyn9I2L4DaExZBbA
gssRRXYI/0CRqxAG9EtPxEwCmf4xuqxH2Z7LsuoGsfVEQO/Cj22VxcsTcmpL6HwK
sRNTFpBp340C+QINCuyyLewijM2sMEzL8Fb9s1heg0F3WXh4+EjWUmiqKUBkSian
ffGRj5rrxaNb3O18wPqXj+BfhKhaGdhw60Gxyc34HJUZcZuWyKSjQmRC8PatUZgm
ybanskts3W5w1Z/O4InffEPWlK5075JH6o35RzJfqi1WH8//QS3OIjaOAqbnbjz3
r08yDbYS1BDwYcDenyPkRvtJg3UmpFNLngu/ppxHIGLpVtONgNw8fPxoqx3FxSMd
B5ic8hfY/9AILu6hiIl4fi+tznsyyousnlKkblBoMCqVZCAB/4HShJmgidmlwVlX
dGczTpksvmvTBDIvGTJwZtIk1eW8B6I9FRpDNzk4OVYvaglSEPJBZ3x+ckC5uvJF
7aXgD8uW5GzT/I/S0M0efAUnGEP3zjDUVY7tWoFLUTUZyQNzZS7UUdbTwe+cb8ix
0EgJeOYbQkrrB+hbIEcUZuud5jqbJWF92ulD9SYC51QlzrRO8YntRkVwK7mdlN4j
OGDLtaneiAuvaPkxu2TSWqntQiDRC2WsmVtGjb4+Qzgwu2Fckrcf1jXn2Yxr1bi7
nII8UF6M22YEdAR/EQByCcTDiMMkaiR6aMxpzKuAvZ8+eiJvG4yrPIgPP8f/foBS
v5Te1bPZ8hsQbZP5+NOtdzn0jafkWcKv5OSzrH76eXWp1A1IwhLd3mqqHMaVBH0k
nAwvtDibt1o142vAT2oR6F4MXO4h8wNcxO3YQc5XkBI6siNCV05H4IEd6CUI7kDU
LSjYhW3d5OEbR/KR7y5eqSQnPfg56U2ccPJALzsngOwFZUXCI3BtdaxDs2560nEI
nTsTmP2xDgYMoH4PRSOW2oOvXtB7kgcv0FHdTtJiF+SHA0rifJueO2SSaJdm/CMH
2DQGDX3LQ4uXkAQmUvsEeIap/1k0hDaD79WebC6ccgHsHY80dH1NKd7skjveSFum
CO+NaHLannX8vHwOkQTTSMcCvBWOXowlmhLKD4/SrNE118K8Sz7QquWPQCtxokui
J+ihiWmw3QYltnmJR7tqkGjgMzVBlXnD/plS5ILUg4JNsVsGJTn8jj70PKJpHf3v
Ve5rDic36VcelT7TktSNL+WitDIonq6Nv7+FKNtqC2TyXV4wdaIWLPmPj5Xk7DCU
+RNYFNmXH6IraiB7W4r0YYqbnuueeTjjABjmkKixtNxoLtNE3cUrs5FT8nVX93kd
R/fX97xuV4LH+AA9wvWQJqWwzHnAP93EeHlSklPXE1r92ExaL7vs/sOGdf1SNgWe
MS51BM8h3MtmGoovkXYNliiqo6ncitZAHLHU/CVUw5rAJxEih6H44sOS7NI6RrsF
QiH7dTwB+IPGLE/Pfy3sx84tJ49ivgjAel6zzVg4L5hakWzQ2KwGBDqdyhG3787u
ddGUJfmQeF2ovnYxam+kisSi+vABp9kOlA1XLuO9F+/FWtbuugM6QIqKFyLpThps
LouRY+eaDFua2hU+pEEOshEEPvdDdzQXl0X5RmDr7tRGTYcRo31n6c5IJGi534hd
pdLCjHHrTNgCv4rx/C0PBn0/V6XyR7eG08MrMEu7xiCaYh84a2rFFkLw5jH9oCdj
TjTwjHtHjvJBApq+UVYRvj5EKUt0gxL7Y/4ZJl2rBzmgUBHdWvPM3QUC5noER7Js
yQohNQ6F7yWeIZG/tXnE+HpufSCxUYuX7DG01F9ID5S5UT8mhLsU83Ml/ezTFepd
nFI+xxhU+ASXt5dIJ3dKk5i87rwnniRFgXrt14WLmSQoe6v14BCkPBT/+0+Y+FE8
1oedBeNGOe8UmkSyxUwL50Hv7Rx4bqrCW1ppY8e5PAZTRj8ysScfJ6NtB4MGl8XE
RXo95edAr9XWUxs4OGxYrKIC1iyFQiyfVjn9lUwERp1iqYAPYZCaz8r3wxMaEjUL
MNLGt5ny/3oVj70BQJcs6IvN20fL7yO96vEwnCwr8b7jVFqv0l8dwhJkFf0KFn05
hyn+HesfnRDY1LJWZSm0WpMqtsOKELLNH2vwEzD4xOoXs47TdPdGzqrmtWhNyeMu
5QWD1vDa78z6iQjGzUumf8zkiPhu7VTbUG8pcOZBi2/TmL4WGwKz1aGQ73LY/wnh
a+5saBGHD2R7M9TBZb6ouDpOZeC0yJerOr7yTBFyex1d6w1XTyGo1kBy7YTsq8c8
SVXHVSm45MWFW+wld4+baIuYOOTImVNLJcV+647+xzNUI3wjJfsKyslxGdd9EfaV
/tNE0ICojMLfTrgwnXIONQHudFT2DlexCh8fdeWJ5/QM1xBjF+HbDSvzRNDkuakh
GZcMJyCNRhkeKSvigExcNrU6hK1if1/JghP9tqsLaDCjAayflRTYQnrjwSWlGjhU
vpM9CrEh6CMcrg7+cgwSJypIp2fhOYaMxuegNq2mgbNhiWri34gPkKCu1OYb5jJm
uqtNdRgYL+7sZJKpgh7pP4AHLiRGH0vz+A6RmThPnD1c6+FeZny4uq+91Vlpv+bX
FwNPFo50BrplQBu4EKR1RlqeeIGkHiSHKVKvsWgDgiuNxtHwPK/N6I33+Lo08zij
0mWdbmOkRfvXdK0POPr7XMDIHvsuytnFpgezpIBHLd0Nz0VPyGfdbLV9X2iBm8vg
ce+QhDCq1TVCu+3l2AP5NLW+/bCmeuUKzRJEv4s7F74jXEedYgA5yEFbN0VkyhY+
+rF0YGR/Vt5TJ23b/607Ws5GNIqE3/WdS+ZNlEDcqCM9Li10yeI6XfiIa/0s1qJ8
v3obmDt3nKXE0r8gmQFxnIBP17Wqy7VATMHy20pZVRPwoYyff9LlHrlb58DXO+H2
kXyf0TOfwzBF+Xp4ZK1V1plRP564bKn99vgXxyoDtpQb3ErY6MBuu8znNesYVfcy
vyZL79V92tONEcMRqP5qQ6MXl0ME0fNUs65/fUG2VAViQ13xoKJD1U/hd2t+g+5C
K0lGu+zWnwT2kTnXXXtqGGyX079IaC/NuIuHO09LmU1bSv3RZe181S3MpAIOX+ph
RW/k1noQU5NKiwC4IxTsEeQL8LUINDTWMZX6vaCcJ0YMU4ZLp6hboyXsNZ117Eui
R3swN6/4Ob/rlFwQ4tY31Qk9GeIv8VWb1eWotcjCg+G1seBA6Oi+k4QVTjCmoVIs
N5AzpnHpyIulhlYrQCucr69egN8RcOsaVbhZx6cwC1s12M+zPb/s92Zg3GKo+mVA
JLlA3+sWBSr4qhpmxRdZjb7IQHQOtqDea+hOAugWeaDwMKew/ewbR2AtCpszCHVt
zHpqcEoS+lPxXo50YHmbZMWDVOLymE5Z45Xk3bY3D2QGrEsUR988QRv166vT8ptY
ZMbVJyCq3vVrfPO67ADWar3Uf3iZrvZ8Gis/VbzmA2KdaibxL2ISf6UB/cv6lfRf
dZx6nCSTLJrGnUMxhjH1WCzKXu1rUOAa4qs3Jqv8ysVmDhKrnQcvJzfK2KdF6CTv
c/ZwJcxnweqpbvPyybOilUnD7pDm1mcjzmnTopmVuZ318eJGXQMWEANHTGHcMQtW
xpcXHyRMpj6T8rpVDx0tzvIe8RtkZQD8Si7HEa+Z96lAq9wA63DzBpk5M4bKXSoD
C1BkzBtqhq42NZh8CY+Z7eH5+ij9TawFaXn/+iXDGpdaQ2A09yaQKKcrKAqtIHB/
mOfuC7Ziy8sZwpJ6LSc80pnrhYrnMqZXrhl8uQesUUWpq7xnW9joiODsUkuavyR7
gF2aeJxvYFfe8wSsYVQuuX7bLZiGgiYkloc8FEPIIiyB1mQWsVUbBbRk9GrF3B5j
r21o8r2NLTVhhILF0sfA5zrzAEf8Wjwztm0R9H0EWzWVufDKYJPHiAIlcKjLxATP
WGyj0LXaSER1A0yBLsgFQm1ayjn/n1FOvcYbohF52MSNZvuloRPj8bHiZb74r9bJ
w8pWUB7tgMLEAW7b8PXHkVd9SnjXMqT3rB2Vm6JIxf6yf6/+FLWu9m+stvXYrl53
X2lN56+Obu8dpVbWKuKiRpTBa7gKZ0EjPyp4bihjmx9Uk9KvFMfLXOIdNl/DCxZd
yxuAwqiaQIi6CnqyHhwhdl6RUpfHP3RF7Tu9hdJUDkqo+SaM0mHfOEcHvH8atBL4
gfrMoRUKrCthUvMSwaLep9YF3sbaR97H3wsXx0R3Qvuq7ipwW6Db+X0oOD4EKEQn
sNFLJgkFD4Wv+gbhi/qKznswIZncwKWny8KyaeZn0rMjMJI91gjZ1I3FncsTnQWo
GeokTh8euX16OAv5iBTIx7IhA6aJSDiwPDbHtN/F+0dVWXT1lCovJXvLY7dlHBPC
rY2Up32IWCmpaH/KA6S2jvfFH+FfN4OHz8JB0CgxIwfV/epdhnWmVbKPm4rfFZpt
ZYtKygJFBxxWl5aI5x2ogDH+C9OugPnoddcN+WV+VaGOndP3sUttcG2ss/shtkWi
SECWRsgRiip6Vcstylmrsap7aUAlQbgaQmZWbZhIpdhy2aV0081Cj1RiWEUpdIKf
9rGqulbwAgVVI56NJXqTMNTOyTiyaD8XySylxxUFCBk/N5l/BjNFiFvqCEZHfIRi
7ttRu6UnownMvyRWuTj3WJVcMXG8JlYN51b54NlYNdFEuXN3NC6DL6rqgRyqG10A
+twO2xIn4ZCJCcn/mvGWsj9V0LcrmsFRA1SpZ+W88NUrWeZVPJ6gOCNcw9bRk60S
D133WVWtBE9UxJlPa8psCY5AECUYwEnKh5DX2c/lHusb0D+tBicUhlhRRAYLGOW5
jisMDTC9N8GYsz3QXRd3MxIAJZC6iMgX2qT5pciP543j9+WJgpABKTlliRNKjjpY
OTn5d0J1Sz4CdIMAQDEdw7lotjKiZuo3AJ2BfLbIq5oX4D8VwbTd+9PCW9Gc+H9s
F6y0bZZS78ONjQ05gflk6gcgAWBoVmac5RKbvKwU8J5BMZutZcPSPA5zNuf/QDFw
+vi0nJbuhieNZEW64RMXz4G5cmC2wDDuYQaGhZIOmEbZruriaLMULyRNpSodqPGm
424wqdTD75uPHrSknATuRmseKD41RBULuuhPfpHBoxntoPpDNWsLbTtv2mgyHBuX
MJnbsQPKL0tyrALd5CzY93zaShynsG/3k3yaE55nuENfOC7hF//YiKQRBdwlogob
AKjA6GCC3gQ2X10cENm5T4c0mP/Pyz6mZgNtm0e1IED3xvF/eA9gSbUxyCjuHVZP
DxbcJdJsh/0P78noJ7eHjxwxkRuxESlTGmtpAhVsU5dTHJVG1RgjSSZ1y0OZwu+C
1ImKeZGswBhGBXX3NoA/kFluDTYqifNri8JfhIu0YHWhot606B8LJuZdDHa1Eheh
2+6iILgxUYIYaeBgF7ygtF/Y+F8lZcOEO2nlvvCeQq1tpiu3j3ekx7ReU8p6lrSv
oZIP8VVQaSBS3sW26onBoOkX8q3nfTmnPmRykczan+LYEwkgMAKW14aeFutYDPV8
/8z2PI8GxWkUi1mUkajA4UGEltfoFaxAj8heWBy4d9FmuBJ/JFBKoGqC/J0JmU4O
Lj6t10WCVtnNkO2FiurCRtc7mAYn0F/VDONNT5yXW8zjTMZX2JNE4W+AKvC8xyRX
ADqTOfIM8okGkPRsq5Bdx8mShEpT+BBuq1b6r5kBCI+oBrZd5WH5dhlelLP4JSxD
fAcR1qc22wySa4ThMi7UZkOHmgb+xWnnvWNE4dQbiSS5aKA3WkCt/YH+c7YLkH4G
dg/UTlfC9OZPeDzLaKworMsp31f4X7u+m4sXg2frzWie106OATnEjuYqkKxuyagu
fctlV9MVnWm1H68w0vejEeo4p9C4IlPWYsd25LuRbVjtIgy7D6OVo12SX9k3nqYx
YuEQVCVIszVws2BhALUEEeaDtUioUd8GdaLntA3g4wcSIid0TIMDk+6v+aZgxwN6
6aOcFQtO8fcvqmylhowpzsK6C1z+Qd86s4dQ3plmZfqU8OcgGTEa4lONVqxG3rET
5Bi4KKYzSHSzmZC/ttR2p+CiXrqyBmIcBCi/klXyhhm48FBeTkReuK+HstzujfJb
wWAe4k0vaCqIoDIbEukFzxWqWHTl3AHJlduDkIqlWi2y8dwyHzsUFc7WA4vpD75R
UDhcCS2KJg9C3wXFv6x4/pVVjupRocsI0tlapsnxfqG7vkLdJzsKKTKEwCzN0gUl
2yCF6YC/ISoinghGy2Lkl4fzonaBCIe84t2nDnYp0aX2bbTPh18BjnNDDUYXyfax
w55AM8KnJytzR0/7V7GHUMejNTsMaXS9lGElvf3HbAwRqONYVV2jvKr6DJ1aLus2
1AfHSsDDOTjNKw7r03BERFEINl9WcQjoWnRXmWf0Ns+CmaO1phFbeZ040DrGVO78
YmPzzKHS/xxIV3wqrFp9NsnSk5SG2F6NrlZ+lAr9sGdpRcdCm1r/Wxwg8cqaloxk
cYT46WiaJada+pWQWI3djiQsrMrwDDdm7f4xB0QhWEmOXfnanM2GvAl71YcRXOD4
apTG8LHeWkm2ULw5Ox58tla+kcgb2GxN6Mu/rTqbOtxypags1LhvWMO2rUAl/Eeq
f/oUmjZy36u/+B00j+QG3Nb/nYPkFXBujgS4l4Ryqvoue+LP75mUmlq0Z5xqsZEX
2SvRcjOObGz9mcxXK7Le4DdmVN+Ab0Zxjnt1KM5O0KdkdoW5FhnaZZ7jR9angjvv
AEayP06j2e+ERM2omvRbhy0v4v4PAMZNv+e7rjdkaZMW3oJnWirfYtIsug9iSWUI
zwr2UBiH0xyUsCR6+RgximY9TLEy5u0HtUcsepz6oXfsDuLwfPCdbYXOOUDTvgBk
jOZKs9y1XKsQrfIMyLjIEVliO0OgIB+Q9Wc0P6JJC8Vao3k6qWjfVUL7I6U0gBSy
n3/iML7VjHr9He4xVEiTLZY9sA3jr13bA4+phsMco3YXySCtR/xrSj4mEM9CpBVg
b/afsXZ+zfaY3ae3QANHQ11lOXRGD8eBLIXK5VEoFTz8iILdIK7GEqB8nALPaQX5
ijarv5zrUNVMtO3wUVAL4GUX4Uddq9sGts8bzPpZDmyaL2q3nBtlQ5gz8tcYrLFe
8593Wf/BgARom5rFwDL02IMmTrfVe0F+CMtxFWDZmXJMqn0hqgyfUvjydtKwNksp
ZdhmOLl/yKcprjbXCfSvstXs/m2LR3zJEX2FJUBdyv715pdwCd/UykNgmTFvVrXd
ieJC1sEbAlTvD59F92ineUyLjKhqpowsIhZ/scjYwNBoX6kFQW3N5nSA6KfAToar
jAUB21CUKtbKmPv9TVPhRpX6MeoT9fMCvT86D3v6yIfYwtsAB63GWrlVZ8+F8qkC
BR62cZrqXLkVGVFxyJf8TqTlc1B+npKF+PKjckSneVRGtP+q/swzpXh43YkBbunr
xo9m1YoO9MnPmktxWusF0z6pFCum0kkXcwjCLFOsAJkDGZ5z3XFKqDAJbn3WKNlP
mw0DhdbLcuYK3mQtMU8/2ZXgJzJi3wp7nC0bXZ+o1QhTLPmA9NS4FkyTK0NpyZ3d
ARY7QDCNzEd7MaXZxvYAT7NEsV9Y6rAZfW/kJNFz4Lvxzxgn6bw3nQTfU1uOPFF4
Vaeqd1PnVBLG6xw4NUZUy9L8kjJ3HbWATkUNJFvdbMvFFLPfZfE+nnQ4MYs1WY9J
s5B3FMhcFr/9Rpa+h/hh/lQWW6HB+QX066GYv0Z0gpalcZdfzNYVSS8ZV4QHIjtb
S6b5H9f+ZMz/8lvKS8EqHNvbjPnZippeKH2mUKLv1GSyFUZd+9sgR2o4tnzJz5gb
zqEszxIdZp4xTyvDYv0bq/KwoGsABKeC8KuLkBdQ4V35sS0bSN7Rmes+VevqH11l
a7PWMowwVXnW7a1yANXTy3Ngx+zbYL0z/weKfPOHEu4X95byyu+np6O+9uap0sIb
XAx63k1YtvUkA9fG6YlyQOkK2CtfzyfrwX8ah3Q2FG76+obb24dgyhGs3yO0tS+Y
EBFxFo2N1GFcx++UrurPutiVJ73Ls0bpAnv3DCevv8ZexW1qgZniaihyS7GNwjvk
KGDwyEl3Vhh4xsV0c2SQ/ErGO27Yb4LIsGTVzN7e6mCcPsVsMZDYJtl0viyVez/c
fNc4uIEYgA3k1iKOYZEsS30GiRQeLA3h3+DUO2h1j1R93cGO5B2beyfCFBOwouUL
QzynrKv7EHQe6Ao5d5ZBRNzRDByd1ZPSUbQSHvCanBe8vM+PTBTilZGYY7y5C9qX
5Ae1+qu1Owgmw/aUjuBjtg7Hot64sBEUSOf4Y7O2oytr0rztNgjj9W9VP0uORlhH
VypZWxLvecoNWOZX72kvtIgAD/iAXcBJsxVfDmUl7CI6YqGal2jUAa60lC6g9Hsa
zu2H+09P+2epHKieAOwyzbvSd/VxMO5AP7Rw57fsUrHct9PJCWhDxVKWSW3y00qC
cta2DlPh7kaEmdM8aHXKfqMIi6oYFHqe0cJjSrYI5C1zapUgv5/c+qjAcvzXs6/x
pVwzDb7FFQUQdCbVYEPJ9ijng1xNIup9Et7a5hbPVFRS1RREd3EYhDui3C/esxSA
9mgE6nciBqY+Q/TIQyyIN4Xc8NKbffv2sbbcX5F9ozavsjLm9ka+NfYDmfnIvEu6
nlxqSphHs2TmjVyoYIZndJ47+naAWrsakV4rK0cJFG3lkkyhPDoa2QuN687NTCiM
6MY6kuqBI//iNyxU+SaTqMsWLCZ1zi+Qv0EMEpP0H6MjQD+zbDtqDgf3yeW0K5Ap
io9WCdnZ4pYSFYs47wMvjawofJbVoXt9Pj42l84dU4UIgBZHS5HrBGse7dnlhYj+
n7V6XRZZDoLpG/LDRwVVLP65botgsGkSO07tmvGKsX2RTJpW5dCWgIuOuZDU/XA0
KGyz+C1cT6g1lLmafuLl2swuzm4iW0xVJ/Qc8W85dOs+XEqshFoQIpLFM8yuhezn
dXEhmxyvBTb5Mu/dwn0R2GDLdJJt3QxojI412xNG9WhJ3Lm/hvOM00eYgKshipTM
96h2hVGZnf2MsTVIInS8KRQu2Nv2bbrRO+6jvcuNvDz3zuMGJmBkgE8XnlLRH2Bk
g5TgPHSWxS9dkCE1zHlhxvaMTLBOa4KnQt4nsNG3B3K4ObtqQhC28ttQAza/uUqK
ovEYPKtSV7TVFIj0ePaijd1dyIBnHFXp8y8zsPc7ncCIGLiLIkTQl2JikE2T/eN0
Q2uFEjxeyKGdsBSlfRY48GL2hoRziV9HGBatg2ek+twx71auhvhtY2KmK2JLQ0a4
DYEp2NYFHx1aSWejjEPoI26GTdoH27pl7FJjZtDe4U+D3ilJXCfm7Jg94ElXke1s
PYZ4sF/5+eE4NKwdyuoOsTaY/+XtDQVi9if2EP9OlwNdcYktzHA5EFGVLGnkVZUZ
RyKVJSCVpE0UV4JJ8KyVxA8tZKZswiXYaT+BNZAOpwlHavqBJFjCNb61FeGgBKo0
pPazwLxbm1+6ng0oTbNYRGQo5ZA5IRCwRtA6r9nhUdB8tzgaIBjYf7SxRUaAPjKk
Yc9Wvm637mTo3gDwEl1q90ahK/NcxwXT1gT7dDyJ6VihgMkSG2+KpyAfjT4EpYDn
q1kET71bhr4mRroctQOUFTfjDvMt7cVvZByTlLDCXxDYB3Dqr/vKJfsoSlMJcihv
eWCjmBi3CZvygPjjOHFy/KabtbrWGJEW2GQf2sUFaV9OB0wJoh6eFrshRmejBOnK
9XOZVjfSFYX0mTjVH2eohaO/6S6FH5o3qTDWKyJyOpHV8kmmMNOs1ZHbQeHD+QKu
X0tKwS5CQH0FBYj19a5jDKKGP3SeheVNVHt6Ek4i94CnHCknhKuItbOfnXj/vPY+
ZUV1DmSzkhCascogvoT2HuCtNuLii13Di/1zB3plOoRgbZjv+tcKgYlVpr/rLpvN
90ZGbl6L4Kmb37AOceLIN5HnMGuknGzwOftkrOXoZpoIBdzl8fm0RelvIVdtQqn2
mA/kDSc0Df8pUk30gy9VOkbJ5BwCMfJWLAyoKEDYKUIjpDiATeDhmrODqDYwcbCY
ovrRRCBxhVEAxV+HPqNM9NgzbuN1WZ2Wew2Ha/Y8IYl7bed1kHYRID33kvGpBool
WH5QwrW0vqN8PJSqT5ARbYOkBTsYZqrdSuCRx2QrW2NDsFtGnr1lWN6hdtHtLavh
5dyYOB6izQDboiONpCUmGz9219vk93EmLTptwxi4CTsMB2bKt4tAScjC03vdKJj5
asGkvP5rkgHOGH8sFNoPOiwcCDILojYTJ204vsc2mVG/z4Oe96SCuK6BVhl2Uzvh
NXRdYmXkU5Vsn3MfRU3BydGH0+PkCkl4hoAF8Vxqk30VoffwZc4TpBrKprefIVj6
5mjEoNtUwyx7V/n3QXmBhcknqS1nNjwS56PLV89oOTLX28P5B4D9cpacpqPSnw2P
DjU4lyvdrOBtNE95/o7hGCn4/+CYi4idSuNEZMXJIQ1nX8V7a49uWxgBC31dcOms
o3AOMZNL0mFdDAODwTtuMuD0qeZJVtKilqJCUkgpkeBgGuDRWpZ0hmj9DZDfhuQm
QQ9VBIsPVObK4ZI1gOmVSoR/0ePQKEIlZiGgZW/lJxY7k95gmcGe0WY5A7AJ0mdS
rpErKYF6QQpbsTy1AgTZrrbrjd57MWu5R5dA4rPRdORjhSoSGVmo0zvstyfoyJ37
AE/MqmoTw+nVZo89vHxwsbEMF5ecdfaGusruiDFptDzFFc4dHrLUrsysh3N2Nxvy
raxcy0r/D5W9YX9Incec3Y9Ks+71UAaTF9G3vI2m0MVDstaYg9tCAAVifmUK3Wpl
EiLQbv+MmN7Oi/qAIrYsjQic0chAsOgiT7jgzLAlxsFiUeZphtwcRww15oLJDOog
rzpu1odgQXuf6zRn6sn6hzrfLsYUI/QMsjK9Aj4Xu6LbyoWPfunHnHMeJh+AJU8Z
P2agkYZhH1b5HLIFN+wLycv/xmauonKvjmBqS2ABNtHwYa2XqBWEc77X6qlEA0iG
4qDRb7wjVQJBlT0aQa6WJm7kpx+JTUECW0cUFSdfuMEXp2E6aaRYrbKvFiGdv8PD
WyNgxegNNFME952nSjynUJmRTVM0Ad61VKI/Zm9RbhGc668XWOHXM7WpCwiNetJB
RxMQ+d9s6b9n9OmLoV169ySwA1whwpD5xAqVt3eOncpQW6Vs02qZQClqvwx8iQWq
PlSw5fHaXoYdmfYkT7OvYoJ0JlMS71ngZtyaiqUq8GXXuG7ta3gWqIxhLhvis8ko
km7Kf4+xbutGw9Nqrrb/GjHsrttPe1Jn6DgtOnQ9DcPYMYb9f0sujLqyqinbNOzb
M11VcmOcxgfzn4zF3us8ZjhsoDMdGzB0p3CEU8tikNpmk/F1cTVe2eLObJi2QYjK
PfMDaghdKHcKRFOEnBziQ//zwS+KdO7K0chTzVBgjUoSCH1+J/tF1NXQ5tv5XsMD
DizE7s2PvVXnkOWhCABPW30st3sUCkNXCIjK8ZVJqFjqoZmLjEr/wP9JZciIJlZ/
mumZ2oXcItqgtJ1zhbbL+h/XI7AZYGbW/oD39ED12BZBdQVS6z3ft05FUWyStlNH
DFO/LesEZzRxHbWgcQSsKbRMzE7D/G1wK2oIUzthVh5RuL0PoDaqVwl+XjCaKQ4H
AHoRBNWGpYAhMah1AdB2h6WaAqeX1WpMQWtSoawdCM7bBQxdq0w7xegdAoL3hdmy
VH0mKgWHZlOgy9AN11QCguFTPWQUZEfHQuSX+7zTywk8JBgqaoS2S52Pd8mucC3Q
B1mx0wl6rH1DPmUXyzmvD6GR8vn0AQbHml+Z5ZBuNdr89Jhy7GDbksH2O/3JsA2w
EH54KzsAIJDzjOmeU7mld36bkoxcIaCrEgBi84F5/pQoOak7Q/vE2ftQt37WQlCY
EmV5diNjSM8DztqqWSIyIQaXjVAFbRuEN368YF7DILI1RyAsq/pp8Q0mxXgMUtKr
5TorD19W8VZVpau2GGFbOMnoqDBhqi7q5OwLp5EJU40p8mcWnkZJQbtIIvXoAK5j
7SBQfT2+QLas/TxpYvfgQFag00cLLYyfEL/n8ebOWK0UVoEIWCyp2uj3jqqA29mH
pHN7hCPxtg5WJcjr+M0O/ioxIAPdDbsTrBxeV7vV/YsL9Zx0mn3t2wNTReKAsQE/
EkAcDD+UedvFywCey6pTE9rWip68VF4ZGCnk1ctJREeFDy5EcJT1iKxbW4jltFAI
Af1WTTT/dOnXDusb3Agb6wSF+mhNfpsAT5AXfFvqe/rR/Gut8wnCi12z6y+tnAKz
9sf/6KcJysEJHLs6uJfX5kWD3U4nPyIixRijfHLNrH4uzye3YnAHMTyvBYGYJGvM
PcRjBjb+KDV5bvXCxTKetDqbtMjP6eezcaIWBCumBUVROZWdOsWLSoUtklqPOA5o
fw56zdgAOuosI3+qak5RWhs5ajNLxG1XFk7lJztF89asztbKokMKkQgsMap42fQ0
MMYpnxEoR+8pnlxFzP8PcTy+/7wc8pQembEbfNw9z5rY1kjCzKWDlnU02es+/PGk
gHhsf0kUqYG2SSRlK20dmwCQZEYaYKhlP3zREkAbDjCcKVXE9XxWb0TsTGJI7rvH
0dkrvYzbF3ljVwXXx6XWpWlzZXXKEffPMDKGkn5XaQ5d7YKONw7R+Xy7I1yPdmCr
Phk4z2rUjf3d2d9LnPHXZtOHKcz0wEA0/4aWW7SLFOIBp/PmvEoQTgWs0fz8uxOi
BNKl3QK+4+f1NWwFm53Gg+A4scXLzz28gAktFd+0lAHq8rZlEBnHZln39j6lwjSV
Qfd6eYAqcOhB1oDYSSuELQVtAfFX8eSZQICGw9awUEXhJJTiQRWKN/3IepmWModH
WpNqefjoQ0kJZ7gdKriGeXwMXyqCp4WN3OF5dnkltPAiS2iH0Cwte9TRivD5+epK
0k2nQDqnuOJ4dNcvo/nCWPqRxwUyynAyLJm2JWlLcEn/PbvRrN8OR9aFLCL583GJ
Z4nREhUE5skHAbmneGUvkeY29nDXYANlwPvI3LwIyPlSlJ600V/vwcBUq+xzCXHe
SbbREjPps2iHNnYMtnqmzkr4kgEDxQAv/f0lC6X8U9FGMdL0JpHYtqDaplwVxgv1
37/IFaNKt5O+M+hqqODthDHQkI/WWmkHDy7RJZOn4bqr1LjSzp2KDvNRmMPwisYo
3k+yMflmSEMn+w3m5pSuMXZ1cf3KaXA/65etlJxtO4UKGo8C9Kx1kQtFBrFjkojd
vIJ9l0zKumTSqjkuG4bZt3LZv5ZqnXAkFq5e5YS64fWYtmoJVEEr+R2komTEZaGD
bjsdO76WWwmAwVel133UQbbgCDDexTQb5tA7FhcLYKKQhzPCOihBtQk9D3BrpGY7
eVQY0fdBBvy7OUeuzsESiduszIk6Itl9NWcFLaeIiaSYQHTZt+5T8X6EzejVN/Vy
9qH9Qv5uc5yEDggzERr78n29FLF606eJG5FQplkksbBExvrkwCz1/yYRuqmo1EIO
FccyQgcKCNQlyS/Zq7MWhgII/xW2cfM/vWrIO3+uhH5uhMHWEkpmR9nPbFDAxZ9X
ObU4jm6AmO3lhI+aNZMlZph3mVkYq3mJe4BNxTF3+4PflL3S5c6NWTe6Vm+QVrVy
qQKWT7M3ecSqURqesveUaSzkv2Qg1QftzZ3IHh5Z0wWjjxK+QLua+kk5OsXWTgHE
zrXKeDowmO1cLrCSR4gWf2k9372YzK2GwSIeA252kr83s6dUSOqmRSaekV2qb1g5
I1rXKW+URhpmjbMRseWNFx7SxDkwu8dM2ElynjWVxpB4mkIdOg3Tx2/VtJ+NHY1m
0StXZYYxYdi77EMXwXHS44D9eKnFizIEI1g4B3B28IGRTr8hEDEASHg+cxhos3rY
A7POcablyBuWIFMn5ZWG4NzC1DMO2r9XtU+JiBLQio0b6GwNo99OCA8mX1RrJJ81
cTKmyVd0gu7BI45bVxnPWb2eGgAD+5BEh2cifS/JfylXBh4iV1Syghns6k4Oc4jE
KlogHVtVvI/w+4nmP7MjH6utemI4J141VUi/8gnwwECzeMCBIRztoJlwwSIloeRI
+9dThvlDAbPfI53vrODS6mhK1nnV5gjcNTwX2Sl7ShJpAOCRp1n7LuW8omXBrW7Z
1gIIagqAmF7IUgLPngI7dUD8Th3tvfgsJveqTTwMcGwkJiDdLQ/Q9egRnDsE9ckp
99uhDejdiK3mF0oklZpeaZw7z6p5JdWwY3jAaM+fQkEBBCw+u+PuqJf61lDkLpnZ
T/Sp7hU2xGH63DMhhzu9Nhv+ZcexEdib4vPTId1eUywA304UGz8b8Ox4BhKnk2ci
yoKAPaqS2MMeljWKqsv7GLFYDLLFNMaOHNeeVQl+vYgpAmISKcffiHPa2O2JACLg
JSYuaHl30sW4uC76AXUUYkhuSMUZEhiNO0RvESoERM7yU0j6bjNgVOeUndObb63X
nHqGdjQ/2S9ajuv+2nG66UIVhS253na2DsxewY7cg8SRJhoQuaEXa/PsFUbmAzjH
00GuATJZ0oJBY+wiEW05hV42AJG1u6pk9IUEatAJfbBr0EMnp5cKKz/r2v52D2M2
t+nGW65z9fyEiHBi+DBoq9/f3V78t2YU8dlFDAlLjQHz2U3YS2/znULyDKeLKO4E
T4omCovuH5welrE+ttchgRhFlqAl6Edd913/4AL667w9qDBeuTYdsOkhHM2wskAv
k8+ZgV5GL58EKmh1HzWoiEx3t3NEw6Zkz0P46eQjbX13JUlLaE37TV0lZVhZl1VS
oSrVZYOmNcTIPknCoPG9ONBt8sNbbevs7co3z0q9keUoffIYJYJAY/aHGp/+3Gsf
BoeZmiUl54iT3a1vEidJGQ+p6EA8CkoCs7S3+3G17pujdVdjBeluCHcKucJdUbM4
P5OhNtCSD7/lz4p/lLWaIlC9qh1eNGNXZyPuerUBh5DoT7NXA9Aj6uP+khzvRUXc
v9fTg1aYJxyOYlzN8C2MLN5CmoCzb3u6qdOaKveuMNDVg7c/QUGSsPk3kED1DIoI
a3AFqzl0d+eNv7MUjTdiDEPQlmfz2iFEq0Ioh7yFSqmGW7WGtNJT28ik4n2PpWER
h9rHHPyd3UP1kpEoXOQrOaQevIk5FB7z5oiX94AZDUDe33tnE0c6d1l+Pq28BtOs
miN3Qg+OO1k5SwaG0Gv2/yqQPGdCVPq4P+12eLGZ64Ilm+HHJoreSVxDlg+SDOy6
R3sg3MPBMYomqhVyTYDpIQthuD9ZxflbDZOphv8eI3RkkK7Ag3PBGXCgRLBAFDRO
mO63aDhELTe27FnE+zy8uOrmshnS68jcvIuVFxkJkG6Q4lvxF2DNIBkIOA62pGvl
dXQyWOsFgOYuXI/FLCMqYZZ1lf74u+w0CW4he4AflIQmKUEcHXkGIvTpNr35xqvr
ggv8AJwNBCZ+q3WxTbaK/v2N2CSBv3XhJRjVroPtSK+dk3sivP0CeF6xUFJexGbD
lR9dY+rCu5ker2ieBWJKnMSe8mFPdi/wpZLF5HdaSQCOnc2YCOOvzrr/Q1vtKtcv
A+GGIpWdzem1JE41+dRxw1+ZoUWIUiWwDyi2ltYZ0F2ggOz6p1nYrBlLNrKstPuv
yukQ2bzo+r/qQaWE6Exmb9hIKicJLlDL1JWyDlPJOwAFNsSKHw5clxF2mBGH7Coe
h1hf/OdMgYJabAOD4iSL6dsmXeCC4VdofVk2Ci/IaD5JDi2fAPEH21OZ0Zk8JkC6
am85qiOjB9uT1N3dZUMOZ5ahCr2EJWAWmLOi6qX6zb+1uyYVSv1SPsnqJus0qmEn
S0iHxKXtBfxUe8htyFP2jfjufUJ3T1e5gtimcQkCBC2HJB1tFlyDSDm3xY/rqLMi
AapOrx5CI0C8KpG1QVeEb3gJoeUx738Y/K70UlJ/2+7beFH2xfrPpRzXX8W8AOSk
NCbesUJQk9BBVJnN6zCv8ANordNWPHxZ+sBn/J/agkVVn8A3BA7KJRYVK36TvSsw
YwQ79WEQwEiohyFpaHNRmbTW/i0vJU3xItwqdO2iectEb3uWOsQPFtaaeBxHkol2
JJqp63PW/OGGvsREsE4zlycz2cOGfoKMw3wMtx7POenfiXEEezPMnKPhyL1sGObk
xZ0RQZk4TbnjgLALjKC03r+LWOrhJoKJR+9GnHTrWYu0p+1sn26Lp70xDrt83FGG
TTE2TZQ4i72b2NvcbarUxkQ2PULpsXMVyo0u1qBxhTwZX80BYUC8/ITnv4EyrKU8
igUkZfSb2+8MOqP4quyJAbKXL8P+cfEv/3vIsNIjoXCAeJniAHJXSNUX0FCxzBSz
Wi6KSYXHdkEp3h7/yr3XrGYNyVjrJkBOmh+n/9YKPIGifzYYQ5xzoCQGZYhzEYRa
iyM90//Wim0nhdUpFO9ES4G4DwNg+TsB/nMaJBe0C8y5Aqy2NQ0Y/sMYiYLnT9gz
6aI5q/BNOYjet1gUpVbkDmKE6P9Xke/kyZbtPc1otFfMl5MnGC+YEm2mQy+Ee7+l
O4qaO9zuUrQ7k668TD5qHytzt3Oj2SnwnlnW0JxLc1dDDyTRCFblWW5uP09KIXS9
unwZ8dYpQWRuqRDWQ4wUuZtEGzl6iCAyu6WOLUpsbpCMUR1hd9svCb3JLdGWEG/H
x1fQ0l1jhVTpXuMaGxq4TMfHSVr+WsZyp/9y0mQSUIDTxSqPmq2KwwkKEkUZBWOe
IxnE7shf7hdeOklheWhBMstM55En+2h7N8PGuvwFhN/GUKw83oXY0SH7sD4mBLO1
M1Rj1tn/4P512e+8c+BPuBVJ/5O3mUHe+SXd10Fr3qerCW+aBM+PPxSRxkKjdM9d
C2eD0kqjXcFGFA5w9SBZTH0TO0QZMDLb5iEtRkqgxTFmljFgNwSg6bVSURnoAUXs
qn+xmPZjuZPJYviXLeqELPfhOHGfM3mcLUnJw94y+tBlMqeNltIgC4okRSUWr/vg
+FcNQeQKuwujUIx/xmMt9un2vLYGWjauZjVRl8FTWVFgGfngefJ3ypRO9YRq7gRI
agRVn5Hr0KRRnckQ9D2y8/VCxqfZNE3298KJ5NT2T/0DfhEP8cJi2i0XzrbQB52r
/QVub/gfWf+FAJvnYHWM0KZ5nXuBsS8Csjb5DXZ71fuOlz6SZm/IJcpefufJvJ6Y
DPO1a/ZNXq1nzA3UhPVpt08jBzg/MiB8zXXJqgr5cgI57bxSYVL0Uo7Y/rjatQRf
F5yWWQ332ATEqF7tKP1nbrYYxi0zfPC0e090R/1ZykH01WCKnjgDg4ipveBCu13U
0PcGQ51Sw6vOD5sKBjuvFAQ1UjebqHjCe96fz4Y/SCNdvKKP+ppF0sJRe1VQw2fc
ZKlZsLMVGZmtcFMDSj8VUc9W6de43LwO7qQtL7pr+urDi9BYeWnGHZlVYagDTzld
q9GeKfzDBPH8JeBFOEWFxgInaVDBFcX3CCjMLdK549KBGUIzZ+0h50HJKKX6gH1o
RDZGVEPZ9GFGnaWNlQnfF2lQPX8/ppB7Cn3Mur40HZPv6UVEYcVrO2/cGrh5tSzX
i9sWKr7vLhIBBLQD70LNNATApukaBIdWaJVCF99fxKG0DO3iF50glcCj+YOfO4tx
4HjlsCcQsiJ++yKIbuABML9iiSZtmeXQ34Oypa2jGY4uj1M/l1W6e3iX7wrRQCKc
MJjsayRXHN+KDMwddYzw3hsiqrYGZUzHWWhu1bZ3Kqg/xPcXxQvvn+FoYAeJ+Gxm
R38zSOo1GY3OXNplP2JbFsqenwB2gR27c8BJSNcyJMmOJNZXLM7PXkiOUllCr3RY
RNWwiT+O5IGvZ/xxDkFRpYOl7IzyoOpq5Favsafw/W8rV5fm5fVDqmOki7+9jYRt
j9TYnj7+oVpLw2x4wH7d/9jYzMd2nlYssXGq7Hf/MMRSy5KPXqsEkdjRwbyZp+gJ
gbbRj/L3JDV+E/2poHCHy6eNSbwi2ILJ+/Rlb4PuvmhT0yUwJp8daKN1LCshHCP3
lFwV89hEC2aQxFD6lbsOsy42ZRYQk1ggcPcCe/auaBE4W8Gcx6LYHOR5Ie7VlF+b
Fid7Juagbuqmk3rkPs4WoFkIgPj8xOpcvymynaVvdkSiIzymVgN/+blF4h2fNr4+
TqubdnvqMAHALND3xV/zdU1hqKQucJxZh4EQP0b4GyJLcV3oQ7VQZRD532ZidzGx
ZtsE/Hkr4VHnDRFnJIj8uZm0EmoHGc9XyTaACioR+0QwsLrEXZluyJllvvjGZehf
PQJ+hPwb+xuYnzk9XlqDz3UERsW8J9WElagJ2DlEyO0uGU14JavAe3OIIBJeoN9G
JXITOq4tffEkWdNjFLMDihu05zr0CJc/3UfRvUiFj61y9jmH5grOX/kUZMo20uGN
2BlacLUkqxjro8UHcfpj7n1mPzsozPA0wMrvIEg8ghptqt0XkP2SLzVMszB/+hH9
L2txdmaHTFPm+JbZeSxUrkmiN2JU3oL4p3DTEQgcv+CTbv6nBSkT2wc+LZpQfnRn
wQdloOX1oNqOpReThL3TX8zF33iZOVZU9SWqsQ8qJSjZOcMOZ9Lz2Fq0SQsh4YdY
MSKNT3S6bxprznn+200hIprSXrgQQ/ZBfBiyCGZnAapgeth4yAqM1RHcrrMNZWWW
pYecUCxLNbkaYcEaJUVM0609ccAp73DHSECsQ95eXYjiAVkW51k94x6owGChbjT/
DQot4MIFhnT7uApAYTjN7UYhOQn6XeBxJIm0NR3P6hkXYZgeVR47n/bOqndbLMop
ZtCj86QqtiIfzOllOP5vL6rPkK+gVHZt8nr2tU3UeLAbYdFRz0NOchdANeiAtLAa
ft1nabWfgoD7wU9FEfBO8plqxlJNgZSF6gOtwvGQaQQIhNhQI+G6mcBLGCFnfFEC
o10CRPI7ifJ6iSQ36alv2kH4Rf/K2wN1FS2xH9Nsa0puaKA1OR5RRbQUKqQW9mzh
VvJPrSq99TWsnXmKy7mm4GuB7zX5yaGWdsMS3QnF5e+ThHSrYo43XVtMvaPKlcT8
LNj4AckcL4VddbLU+sfgzWwfYzARNwbTyGkICl255MaTdfL16KX+AU9AEWXusqKC
McuGC9QYC0i/wPYj3bWg2GI5hB2HXfE41oq1Ee5hHqBvu5d5TKDmRiV5TeLih0aP
n/H8EQH311T9v5ONZn2Mqc660ihw/h40a8MC9MangzzJoHkeCSrxPLZi92c4zape
QMzxxVmzaPzmobWHoyw0Tb4FDLHgNJmTA0z1kIvffwhoKL1P28HeX3SdOF8sqrzj
NTHCS/2idIq1l8VQYcQo/T6kCRRrYzpmX1jVOwcc/l179Ue5SRIWGLvv/el1l8Gm
ZvK1qkNb3KQilV3TSTTnijbqvclPS4rSsxQd6vxV52HBcuimga9CJDGFGGJoSPt1
3NN83RalURpUMv6EDnPMJ5LgE4FDIH8aHu+cybje+YEphOuPqEhsdSxvLNbjw5BJ
8KNyB+ssbaP82pb2M6ivyAuOwT40ms1VNkPGFVQ/IhfbbwmEZg4ZF9WP60REcLPL
2tNLmwgO/DFLaelJrtv5TtU+6maWFmdqfXTRTMCPsMkfbKL/p13pIwaXD6Wb3ywi
ZfDd4wY7i9vftOIwClCnYxRZbiDGym0Cms1M6t4M7Sv2PmkXPmtsWV+NZdtmQylS
A661Rz0sbRSXwyEFXsVc7SqWd0/CcTt0jqcK2KyquvqAPe0sJlBD1sSUd92tm8Ph
mkK0eBiSaOOzsbbKJJ0wWrCw2pZRZ5fn4jXB2f3r9+CGKNeuS0FIteWhv9mHjiHM
rXr6KwxzaLPi80E+dELkUwr++hE3nBIlUK4GTb9HLk3q/1jOalerAtO1Gh3GYc1i
HjHRtkklWvqUvjj1XCaWRhmrQstuDKiwMSAY7eIGN+60OvuNMN7gUePZmZApxG3G
u8Im6RcYpFajdEDLP5Y2/zfgeB5vNuhi/LovOPVqyABiJgn5WcYYVgDnChzY7+R6
a6fw8bfGuX6bZErZ89ZqzLbR69DkecM4FTfazYV4+s3wd9UiYYN2pL7v1oZn+Hlj
llpixXBCOm0Cs6HXoMqauhsVwGjWJ0wzDkbKdG9/u2/16Jo33IwM/HlnVhg3SeQm
pSdjAqLji6sMHAMusBPJodvBMS2fa/9bXPyZ1PqQSq1pLm1IaW20D6oIH6sGKYYM
s9mSzVR1dR6QfYEc78d0Pe5vQwGFhUFxe9eTjJUDtPyE8W8aydP9/XrtyqJxyM6U
j54BqmHl82kOyOLKB+JgnQG9VWIHrv3eRt4aizxNCp1DhgyerNMgv8moju2v55Hd
JDTKn0R/XnnWi3sw7UwcS6+SDAqWgwk2Gyp/2AviIKKRF7qNjj0xPNEkaMyKnQBM
NX0mWm8v8OeFZe+Q5Gjtfcsb0qZs3bad88BI/ECVB2oXri7eS0ZoAtQ2qKsxk1H8
3/O2wakM6ZJ/eBGDB66pz+HRQet/0Maj+s80amT2hCH79zZvk7Nq+N3sjrhAvwwU
SDNLjorx2GAGqpQkdFqeVH/LaHdLFLMkNbQOl0eirH5Pt/+LpzjvXr+g6wrwzRDm
fC0X9/L0l6m1F3QjcM8z8YaSxfl4XX/9+uxFJiLHSlgyTfyLfY9IFDfHJ2xEjVNJ
A/7ue4i5dKeyQ07InvoybPIL0y04BxBPHtjOedvK0uCCuJcMiVtbXfU1b/bQkyOI
XizEB2aSZhpPNeZr3w4nvMaFBPRfY2xBjXbvyLeFOthea9J3kSNtQT6RQrJ43qCJ
xMP8B+NGcdCd3Ee/O2MZm2ZjP4hMw/WxqktO951NRjD7C+NtMigYSzCfzghvORZC
AT8XaDcbepEU5BK57fATASpeerrByIuVm8SWEt3cSkhbBWhteVoePAlxMpb/v07r
kFkKteCfgJRbaXuftcmYWzndV8wj8uM8ggzF0pvu+NuEoelNFgRSxwGvwFCFy94W
8Ox42x1HohlqMd/mIcG9YBs1MNsgZhyXoUNq0eCVef6T4lo9CgOAOvYWogpeIfR4
LpyPsRQP/hmsqQmnoki2GCpxbs7/uC4qlD/gM1StZ1Ezin550Np9qt0czuBtsMRU
iJo3lzyMsTAOmnFf51SeNiA09Lb0jd/ehFJCkX5UljTCr9lNF0YazJURJd28FdnB
/Od7GAfnzf3MfDL3H774uETk0iFZ2+dYIixliNWBxZY7pdBdGvdmNAr8+ZoY7kxd
SuLYIjWgDWUG0ct5wtshqvakLYDdnNOI8QLo05/fp8Zk0Sn9ZqYhQNQ+tCu9oEkm
Apct7XSrELmuFdQtMDeJ8qxp9IJz6Dd1Np4xxJAx5QzFM9OjTWqUzYarCUpFjFuD
qsjJB3JNVRNJ1/5sG8I8O93TxKFF4gibmE5/B+2qD39NBRqXuAuahsCrdmJC2DuM
6MS7d51wSz39H1WU4Iuq4lZVs2UWB9QLnp7GCzhGAoUt9R8V6JqiuPZUJ9w1dkQ2
5Y5ZCJ3FPvcXD5oQHx5USzltRrw+J6DU9vTgBEMZdCKOi45D84o6iDeL+poNv/Bl
o4HuFYypZSfR/fD/bg2yMU7dxekVl4YrVO+qZ2dVBQ4s7IzJIo+p3a19D8ZffjDY
nM/l2j0LidBmR8sVscSYiKXUGL2B8937Uah5TzLeTRY94O+MPGlIx4xGpdhx9O23
+jYWj/y0A3O3dvTU+FJEGSxRmUx80J19kmR++8iGv3lHQz9oME9qeOSpE5ktvtEs
VCH1cUUslaLBBoc7hHhhpBEHAP0zdoKlSWckUjPJohn0SqKCCigzXW+SXIrpjw/z
QxEz/2nklAFrl0xUD8gKkSYk5N26zeXh+bu5MwscgUtYYwRnTlssJpL8EVURNhI+
9m4KhWLIfK0H0XMsuydOY4JLyGE4FVygPT1Fre6rC4Xe0JCw9UTVVgfWP8hr7e8s
9IQ+1U33f6kYKZKWK4b0fg/Xwzn3xMD7EGH7UYfIFQWZbNaeV7ZWjQ3T2+xiBmBu
BkOUwVe5wY+RxpaYizNjRn9UEHa7j314QemTQAA+wpBljerTXI5IxsPu76TmAzsA
1hFqSbiW+GrIwbx4LYY3H2Y/fDqa3/g7qeJf8+pyIskvNCszC1pb5t5IDr90IWn1
SsCDYwymW6xvPhRBC//jdJWUMUKcGjFeLJzSnwbLwTaqJLNdvttn6DpkKjqVXeQC
i9Q+QaPZRtxnqakifTHP0aWyHO97VbDpCr3QBdYhdQkIaXWgUJ0UHCJGeZRxctbC
Jpfu8J2b9xDlo0wX5VMEgYgAkBjq21sCy3mO9Ez4h8MN3Sfzop8mUSceGlM+rRbn
hJddU5R0i0UXeycEACsx2JSjhcKCEkmRRpzT2a8PIXqM/eRCDp9hViw9orIy3d8a
Om8G5L8dZH9usLxxX92fSrvO/2uwnFhrwAx4kK5qgw56JDU+aW3p6tc1Kil1PZls
ynRtWIdHn5ZReHYsL+5mVoKlS5/gJVapBhtKl04t020SNMwV5WROGOPpVm2lg6cW
drb4TkNBAn8fH2Hf0M7KaX/9Og1MxJSc2MOUruIik6SzpfdbZbf4Oqm4SYoFtBXf
Kdwdmltb2Q9jOAlnJUZw2gL1ENS0zfy1ntpCMZ2AvVDQ1Fb4Xv+4QF3G5zYXqS12
vZrkOMrsTg4f6HNxDVmss/5hCFQa3H9trnQRaoAnCLnCL1gOMo0fZfU/VhZ8NdVI
QIrOfV9/TxsteCPqRa39D1nqD8pG368pUvbsJeKB4NUo8yOYNMX2loHnDyj4ipzh
RfD8NM/ymjgATdbHaQB/m/CEmlRmbuiAG88G0iD/DC05GGH4lQAGeiY7tHUuIaUa
+Z3TQEryneq07vqnxKwz2l1XLGjfnkG11X9fRXeAtNZ1luHRPLV+oUL/1hFAPj1r
2WZaVy/nCiBdZqSFD6mTqGrpqkPf2aQVeSeBF5RKAswdMH0tnTNX1Gqf7TqDlcgU
p3IjwrlovZyO70dZcfuFKiDHfO+rd0iKsX6i7oH58zSSL+XwEAmHijaW4SygGq+B
3DuMjz3NnurHyNjvlLD8rA8NUCNZURy59mpHPtyzLSaXb+aJpqFIgB27pcdRcYHJ
DV1qwB7sTOBFAnh1mrhJE5d8wuisa36tOvQrAAL5xDJENPwCv0KAEg/5SAe1v9RM
DbXop7ijBTzwQq9jWANkVkvvhC5uGW5uwJLA6mxHuZQnK9Mq/0xGWKt+odKsR281
Kkn40YUxtbfm/jefxTLzrDvzH9to81D9Sja4F2GPlzySFxsFq2fZnQfoVjEAGeHh
3szG7TkIURJO9gdyw6VUPQ53flTj6eprChuF9bVY8/rXlomoPtlE6tf2Tv8Lx2Vz
bRCo/a43JGqQlK3LPYfYxbnEzQkVxaFyL3xQJiXgYkOJNRU8lfvQCsPBPNN78a3q
B0lBiEGuhzKts09+OYivrmZZlP5rcBo+UOU4Ul6ndQEfLoqWXPEQbzR5/0ncITQX
i9M6Pfjv32iSGWcgWYbEO+GB7iJNKr3WHYNnGHOXFlSHejKQQ7L2AA7xIS/B+y6j
4+OX6Dr8k5tkIhPnY9Mw2sOrZU4Hz55f2KRprphQtbBVwdlRizAMcKOO7KOX2ROf
UTV1Nn5stcu5Xayold1T9bl7yAwG/K/HArWNCMR4+d+TXMpUZ2ioIcy14n6h0Iko
g0Xo2JhCCmQ5CFYiPaoJ8WK4LPRn0yr49AQ0jH0vntEiwLzx4JiyhhKZeXzE6KdC
zc605t+iFfa4Ug2/bhMqoWcJo7y5Bq44XYGMv+ZrrMkPpDgXrkf8jxFbSZjpI8xe
YPDV6oUVgw/U2ZNzGCwY5lxQDkSnws13w5r8kwQ+6jF8DsY65RUDc/2U6UY7OmVf
Ro1O1oi2LxpM/KU8Zg/3o6f1B1GeRcwXcAPEIMtkeBOskN/eTBW+D6vsosFmENv0
EUrENwvev5C/GNKPiYYozYG2Eu7Lx8WbVQcyRqaJbovH9q7B2JMO5CO3cUgzGWA4
OKqCjbol9kru+puiO9J0yrr3z20gidJ4bNl5HZczOJu6NEk5kXz/p47bqHsnvrzL
kdABjeyYYIDOLZzE0m1Biwz1i8xX+3Lewn+Hty0QyKTG+7aXrMhACiNKWBLL5WdI
XxOzMN7tk6rQrTq8TyBlJqwzW6KNsPRsfjmle9OP91vPmtgKnjdbizi3R/qrgeFe
m0jl0XceBGlM1tioOALwTLpDJDkjzA4Me5obXOBFLKWi+t87kbvlgwSVRrizoVAT
GwQ4Q07HB48gMZtOp+LNRJrA4i/vUa/nLEAABCHcB7GQDA0Ol+TZL99ZizuGg9CL
ikmlVd5JU1sOgWCv9bPaHmf7S28xeHtQlcdU+6fZ3BI4fNmEvdYbylOKZTzeE4Mo
VY8GTyxzqw5GL5IOVtRR9Xovaam44BggaTt1YIqzBGKMC2g+l+RJpMEGKj1djr0U
qPz3Pe1XGobFuqNFF7JEGLrR9rvQdXL/AoiTQz3EYAdUKryIOgDoS1iYOvim2SHW
UX4gPuQTR8SF1YOPde8FRNs+7MnGrytfmi53qqXVuQZNohDHEdBObhLKqqVI9gbY
4DqUGiNMcZv1L0Y3qnsr2fEbGn4ConRtmzwGOVEp92wY8ifqLMyIQ2prDEoOkx68
In6w/+aKWfHlxyQovK2XT4rHpKWLoXymBmBjIlX5ax5epoO3SBriwcEMGyNCZI6Q
2rINlzGti7yVGY/EtKVqWlR0y2SLJtnnchozyjS8iMHr1AAWkpRZkxjEtF7tURLu
qnlTjyES19pwaYztX+PIL0yRl9NAm0rBLJIyop8lKUoYQFnbOsXEyikoc7+DicY9
rAKesb6Ip9FIa/iioIwhZG0He6QTmL9dX7hPpsmYpOvWqhYPxZK0Jr3clWVx269+
0RPYgS5RPyFJuBg2IfjMnjM1ynIyIbARPhr8Ynjdwu4PRKN4sgy2POzPTLugguzM
SVuvODRsM/YNXhGaVQ6YXXziVXnBV7pFZqZhcnc5g3Vjr73Oi9P2ZIvku1KWeps0
+Oqd5/lT0XASpLOkZ/1/KFsFjxAusd7fupFgRpTVTYtasoDN+pN6rOhJgerBYw0I
iV6XFcFjLI/87RKBnpjfmCxeTjbYe7+ww84aUb88ytb992E+RLrnewHYKcl6Fya2
sef6DqtCp6XnAwJtdyRljPf9HX6Z827/x4QZ9A21MbNGSXEurlnWTc0jcvuPHMC2
6SziLfQ+oS5L1sAiV6iCURJZrZrM/HlWYMF1h8Rk0wtzCqcxaCyMC0PnaBnhA3wK
9YJvNoeWPhrZkusgPhTsgI67L4WS1hBeRhmS57H4eHwrDtu+rB242UlXyWzMkcE8
crvk/JwIczwbjhRfIzJTW2ygVIDyiOkgFcF6yjDeUxkLB5biwXSRxXRepO0YOgW5
LKJGQg7GNMkmpYdEyC6rrEYvWWx7HzigeSX6aFM4gmXMVZ0xJIEWwcqil+fejHfR
8kcscnBZuYPo8A2/iUeAalBy0665OWI8a07SVLvvPGhEXjK+cXbCpTl0Bc8vduhk
75IN6RbANMu3ctwCqXg6+WZg6PYu2lfqWZzKW4UgosVDwRlCisqWjXWVJojFqBYI
BxwgOxUIuZZUDa0gDgAc7duKY2d2s0qjkphK+OeI2JaNsQDJPxXh/BHy3EsH4lGj
U1D2kP7ebak1myrnHQI9A0yk+IHzSX7XYki/P2IDigKkuGIR6Z8Eo5XdkZE7tH7y
Pt3UTl0It0mgnk+tT9tOv/D8osvvm+nTIPy0fQgWNYcHIaYBpVVVimzGSD5eSEps
6YnircaQKDwl2FO+woHKK1UCvPs4Uhxe2MGn2Wf98n1KfEv3wLBVkwdKE1YTYet/
NjHF6yb5xpudDne1EOG2TKDT45Rm14320FgLyFwMfASFlV/e0LKm32fBOVroN6h7
KdNyoaxb5rmZh8c7mfZMnJF/MK31RezCcQ7oljmPNiXa0CWqb8YNdOGUL0yUL2vh
gopTQNkQDpS0YoyjhxNe1MGmzjHgT/hMX9LNGqP9+omSBmLZDrZTgFndQgm8otm0
qqcWEs9gEZjWWF8lZNm1yiVyadKpQp1juo0O5NVIXtZ28M56nN7HcL3jhvTQHZbS
vQsJysDYwZZswLf4l1fUgj81AmeEp5TiB5HIj7Bq2NNjdbU+C6pYPAIPSJuZ56k6
fvWbjFNdtkYfBjv8a0PUvEC+DatYbcqnD2fh8ZKXRxE62JwLX2UYowknc3uANp5n
PMm+Xn6OKScTPVTL7GMXWV7r0Z7dfAvNx9AUjqvOi7DLJRfYHCT9niAVlDEnamsr
ZVlr1LiJnt0vzABrnL7OLN5rW5+WYI39pHQbB4lgGNlV4xyUXQy1cQXgUPtUkFai
yfhvQAstfkd68AH2JD8GYSi5MAzTZAvLszuVYW+jRjQVX4PpFFDocNejKuVXBcAt
GXBNog+Pubb07HfRw3UPt2puZx/tGkIPEsh8sIrb9+QbtAFUBEAhuIXfrVZzCHNU
PMn3/Su9gdcHAW1YHRfL+SCnQe4v03p9mbI6eZcer9Uka84U9freTbsKj0CLzjLe
CL8w+IhksGA0hC5bDDYHFehlA97O6ZAIfGtBaL/JJQEM1jGFKn5JxpFukbfIQTO8
jw10LuFptbPyaXbmqmtC3u9+9XPzIeL4SsS3bpbfV/DwLEGR1CyGaBzMQnuOWfQ2
iCTh88fm75J7PTcP8hB5w5vavJooaK7yaBUyCFFfG+319fVV66OX2XrtzkVG48WO
K0uQXL/lTD9zolz58ei+fW/OaCGdZmdg9Yj3YK5xHltpdmnRUa2wHWWExnef1BBi
d/N7YT6/l9sVmVYonbc3TX8aDnxckhQJPa/qyg7aToZ9TCpFBiNd9FUNjfYMQb7w
DlB0XYn0WSXX86HfjztVSJdUEB3Nl6chbkBwBvXOQq8C3vH1Mh/rh4xjC8byARUk
BamYP/AYddaEFWk7eNs3+hgOAwDfAF0CGjVq0IiVWTFsW1BIFFMhJVuuex6iwipO
4XcLYvx/Bha4d4uPU5EyU5qGa4uHDnP7QI3VxC3mtmKqXO5V4ewlBwriFmvmrNGn
llUA2wAMPDOtVqjh9RwgH/AwrpHPiLhwNzYAuVEUiU15Rn1gaWNNlAxIQb95D331
e4YAeQGtMeeWT/ZohkBZ7ApTyjTNr49PbqwsTnIvNpBqH3tGiBfj7FWygKcHbxUY
Hq9kY9FoP76URdp5T5tzbHzmlIg+mMPwIyIyJ6+Sj+2wURNSRL8RCV6gMF0urpbd
O8SGps+KLg51jVc5wTHm7NVMzQbyNs76UWBLSDI1+9bnvg4ybanPZ7+ExOl+j2KZ
svpbquHlFuY/sKiD0NUe0xCROsZiUKeIVW8622tN+fj+CmyfT85ceXBfFm5agt0q
gADQ7CV8s4Uo3rXd6I4EJe+i1VVhlLLsimeQCTcVbZQezLzMQfItDze2MJy1jLaY
xff9TWqnuSjkLM3DEdEQyI2EeLopI4T6/WilTqphEhdznnmDDQcQXjoHhx4kw0aT
0frzxBkE+dpQLJReOx8NgwPNx2FQsnw3mFNjFChExH7nM/5lqW+hEUjQn0V8Fdjw
rs1Wye4fOJg1vrunFesGFfLWbwi/dwD+404y9y+vivf5qkfUXjnB++ScnKbrEYJq
a/oC4pZK6kDehGKxR7VNwfetH3gd4nTbtVIwnQPmgeg9nN0U8+sWKXVxefESo2wt
yIZdzq3Adlb5QnClQ6hulweVcSupln20e2rHr+pjwTNwH2PCtLSxAyzPh74OQIDV
tFURvjIuXCbc9912TH7Fim3Tcs5ccbjOrNWXyLX05xhX22GjVc3xeJXpb1Pg8EO8
zXZs3ELmqAdmGrXEL4m6ALCEXFLQxB2OB+ML0uqCPKmUCICiOfPd+KdP0gHkrfno
zqCB96cllp30EJV9GYXbKJU1VGLBIi/oss0BNa0JQaJVR8XVmVbpOaTv8XMrhhwn
BSVKQ+nn6H6L+ch/5QyulbhX9Cb+nnGw2usb7hM134E0VT/nErOTGKbL+8ZpiL4Y
fMns2eNRDSHQbvDniwNd1JCoZnsnB/cBkO9D5sCe4TUFn9vmWGOpZDVXpsCQKhxg
RMUHv0eLS92rVF9RhKuQL4QqD+/DZmyvHn/RbSEGMIK5RfuM8Wr1vYG3m9fgMIl6
QRniaYBYDloVGqYXsBpRM4KyA1O8qBXmDLSq00k9dtg0KQyl8tWZcL+ZPdxObqfL
ZvfTvKmReZ4YLx/SzqV9iij8vAqOabr/PRRPk3pQ+UJh1nd6yhjbqnWT3RwB9Lh0
GsoDlAIqe2xrVyPcuxqbjIlF+faudeB5AL/lUyYmzrj7Ul/bqmLvo2cy71LYshJo
n5frZZEIGfkO8obRBm3Fb6QvvQ05yRtQI/4imsT16XsPx/34OSqAwICIATGX87UC
u2JEY0OUcOS/o8f25ZlKve6RopGgrl+KWyJt5KHHlPtFMSC53s8B0kOq7TqfuBiT
BkJiJTsPEBSR2caRERnLHxcLpdBfNIL7VGJL7kTF2oo9/ko7X90TjCjW2SFLZR9J
DUx+tYKYVx/5gJ4jmRjSIqESaVfiuhJUmr/wjafGMTAxATuEIAE1sbHV5EA/CJWH
BP/iN6suA8KRjJuUE6Qr0eCEeiBeLGru6ZP4dgB5t0CspagtXuDefP1R9WJJel5K
lE0Csb94CSUkpHeGGgHvCgC+pBMXSwN9SW/HL3Si2kMUoeV+Q+qCiWXvifW14w0n
f0/ynYUKIRnhpzkXGcUPECmZT2pG7cQFQhu93hICW3L9OAC9BCKTnzqAgYfPgLqJ
YqVDuRFuUYvujYWCZSFgeHehVkXg6dN9SFDe4cQp9YudYTi32i9Q+dRxwN7/j5kt
/K+bMuITNDt7pU0Qo3SR0tWCUwRw8gV4VDSEO3lD8KZ4hPJxP+LLD/2T5lCgPZA8
YBBOFmMBqpqp8LrSeUVemag02ZLSg4/AuHG6efjqSkEtfYFbvKXCYUHa7u4Yw2QP
fnHbKFCjtFVg3Ybzz9U5yCcBCjHlkwDqoydc+Txl1z4/xSpyCk7jBIg74yScTcij
kiCSGoHzljAFMX5QAgWMRMahJB/uthdBhNol0Mp41wqp6GpIU8xgeS9nm6X4P8z6
W4QlX0VXBEN2yponeWsC/FKb9Kjcy8lZMRu5JLHKJIfKl0r8pvRFnUi/h2A4tRcv
QV+3O20gNGmCxQd47MmyvGKB1W5QCNTrXZB8Foy+/1Trw6jB1Q4JZ8V1WAk+wcFa
85lQDUTxI3BsQa7sLptHdaMaRKcDVDSbsDJvQbzssL9RgAnM7uJXSdDGko9rnAZQ
hjftKtFVRsZ9va7f8NVCyg3VVHSqFvNNagcjjJNIGem4OijWw0nbrta9VY4fVFR2
9KgfKO5DjG5jgd4cWlwXE2ldTB3Bq8qTqTB3uqSC1ojd2tCAR8hF01RKiTiiTYpE
IaZFcx01wTov+YL5Vjj3OOPJrODGgNbkZi6oBnIx8rpZhcY6sGPNRFNlgXN9qEUz
VYiWkBJjVDa7TC5hcgRl/PkUqz34T9bP3U5sDimODl75ihd06DxFp8vP8HeHmz7i
Iyj+mxhSR3ZNvBiM9rr0uLdRiATn5h4QLg94A2CcGyoYG50lV60qdLgtuiKa97LL
m/+fKrwPThBMcD9G+z7ZeFqejZfSFQy8gN4yy9SFsqDIs9Zz44ygNUUxN2nRjISQ
mZb80mlvC4qBPapxkvlFoLz1q9hNdL/3vsrPWn77QyETmwlYf71IXd1ADWiXvYBe
/dGkMKCbNDnCQDWNv6fZI92GlhB5KptfR6JoezIfRMhzr1VdPjFzPMSmhCkX6iM6
ZmwFiROjKyzkGVA8M3ZabVNVodqKY/ibWkho+ygMv4TxXEQkUAUKLkhIaYrXQTbu
jRjTJuiQodjqkNwGih0+3JVR6J4KwKGeqrU7PUkSaFT7DXSntLoDLUxCwuajiAkl
bi4tjoyGHzrgdMXIHNt5jmKyZ8f755oz8jZNR5NywQTxVihs8M7fb69b21ApiSSN
CL3SjuLaweNdtOyBwvWRY+C+2Kci2bT6qJzWS3K7WUjeJrrcz9RUBm0Ib/OQDrfU
tpqhj85HKYnW/wpkNl+EjqIAINVud37RDQ+C+ZsBE8I4yvQkxaWYNdAMSvjZO6j1
8ii4dARl+K7tBgxBI7IzS2O7wPexxLQy/Gl8ZMKh9wovGRmMF4UxBTdaxe0ZnHnb
yY2hFLIpWW9BGlnLurFDcL4ByRFYo55lloXqeLRTBU9yEshkSF/ygaoYhLeKnTib
az7UQTCbjt2tTkwZBIrF6oH6Kceu48AcWQBrUzKHXjV4ocAO+Vn2jQp6Y0BLMBtG
bvtZVpSAQ2/X9FgirXdi65uHdUpZTnpp88+CS+RV8hVuTH6OOxO4WQYzBvqmgOHp
iVK7S9GdZHu2zkngd3ZE8BHK4FY3I9a1enZrdKootpXmiODtcz7d82qAYLUjJXhT
cq2EaHUq8M7BjEr+rM8KXBylu/bmm5jiNp2hw6N5k9NOvI7TK1yZ/cIL43zpYStH
WP0KL+GOONya5INy4TLKrNP2Ca02F+reezGg9JCFItOh6pC1hKxYXEbmKj1JnD4f
kGkx+bTAtkz+lpwQ8csQcDZPRWPRTdi/pbC7W9ip9vvrJyUA/ECfLge9JrN9w7ff
mfsxROgM3SpK6kmDs8ezd75WoVi+0ylNYC4Jc7+fYW3WdIRRED2Dw/Yc3cEUqa0S
FOXk1ewwvW1gNd27yLO549+cRW6j3znknt8L0w9nEXee6M3ci5Mk9RjDiDD67ej5
eIF21wM9Cvd83DXwzXYj2bnEg4of+D8FumvD/kqxuthti1LvIL+mJUYSf6Jh2LH3
JEWASYtJhm+62WDlbcyB/r+eS+moo0BSeKjbBzrKSvJdAxmOPw3gppi8KScr/wQf
Sofsm1rAedGCR6e8rKB4Q8kW32v0k1I4KcC92lLTGhAPDWz+3v6cSZjLBP4iUvO4
zRITS26y/mfa7gC0+GLfZdODdRJ6S4x3smuLUiVAynPU9MKMrDCXXe1vMJaJ73c9
Q8eMiimaDzGN3g+KB+0fRengLKnfMi95oGdA6nsWOdp/F6ejTilsMAeAmBDa0u71
/iyAM5OjUFXGwWtjz3PpX3noIMnILSRCpINSjg+D4ERA2hOg5SxxdE4DjU+GeXW1
zuWjf1aCMa6NJSt9bTs1LqlQ5YP5GwyZdz/YB6KMNs0RerPOMMd9yEzLFuu88tcD
E0enx3QOYmdYVEorkftAWSUi8+Gk0PfCuQ/jr6ygsbafDAqB7S5+dVKIceJDZSH7
VikgmjCrEp/2OwV4pNbuz3B/ksiehRHm+8VomkEr/XWvllWgbcxxckgwsANJ870E
1BNd5okjySrN+iDgtUuHiEwR3bgyG26fIuuQGwDpwNEXUwRFCaR8r6VXR2ZHh9IT
GV9iXvXkzIb+jB3ge/D/p6/zVVLZr3M1Zim2UK5I93ze9nWF1iovlAEKJtqsfdDF
bqj3hyDFbWu8v486cjubK8CRtqZwpb6q0hz9mFT0aeQRCG86P2dkmSGFTEznH8vS
850qqqSmIjG0s2KA8kAqBKwlDy/cOFMieYq4w3+GceOf4Fjhu+5usYCDA8/PB+y4
LvEbIqrAvTbfn0PqViLL5w30uABYJbIS+KrMjRiCZLQQK63qjQDABQ5ZS2qWJSQ6
kgvQGUdk67XXGc187y4129yyT2iBJcZ2Ne1JAko8h3rdKIx5JaSR+bs35fpvKCgs
GrW9LdMHYvDU2e5tPCO9Lo7VIlQo4JHC/d/Chdl1kdQGqNX1z7jYL4onlGP5zQJI
tnwp+lD42aMXQrNt5/swm1LxoCpgpw3/+CpqBKZ3ULDbsb82A8QTnQF1v3VvffnU
SkUQ33Qkj+BNGiZJb8CHYlB4LEfBfCvVjMbXPqGoqVlMG9PjW8zx9zQtvskEQWAy
vJSu0e/m2NQBls6V7tHnAIkx8ITHNG3E1GkIEofOEuayMeQ6IXpQ0mEqJHqwY0Us
o4gb0hshrVsgcnqTLLKl4J07SU03Oj3jneC3qvn7NtArB2/yk3hw2/gCpTXe6RhJ
DtpmV9NLuT0fbFiBuytduEcaQD8Yq0Nwimq7bgqUsYnmzAICIKGmL1dpZOugI29q
io476jDAb4GY/SqwDhQLEnzbXCskYWpvqQVdFyz2GUe7pTynKXkFXL5T2jwOlu5i
VSG8xQVPSXkbYrWrYPjEcq7WLFjd31Q88E3KlSfNWE4vsSZ9Wc/UULsxJ9SDKkAq
id5T7PRRhdcxuKsaIeNWsoWincbw+AytbVBh+edxTKXH1+4xJkE2T0cq1LJCGhLk
qR1xWCNoUwOiSezbCycVR9a/kDWpz+OLcHZDFL8nMOQBdWwKBdAyLk/TsWXpZlVD
Daukx2SCpYLvzg9M6rA/1OwkDxbuI/nFRlLkGgwNAlnXnCRqNuiucIREpUisgfmT
/5hW+lT2XRRZ/fnt5PsulLg9eZqvadLOTdpZjxv+mjdO7aM7btDEwt07/UMrwgRZ
ca2CjErJ39eYZGyfBzpniqYFwqfsB3PwCdbTR9ZegDoV45Aq2w3l41+fURw/raSA
Z3Bkf2IfnDUVymcfjcbJH90VzgcQXUkFuudUOtajP/mk9coRHxsuYkGs0ZgQ6bBo
shqJ5x3aL96jpQeKB3plF6wjtfvi2/352tgZdxpg92vrcPL9B1jAh0YCcLImRC78
EPet0zO8MqQb5BqauotP4wfoT35V8pxVIOEwOKwASwRj0SDIM0pcTrFJD/jySK7s
J2BIp83bIKZWnmR5fqwAZSjaMvR6azpifbnCGZaEFwS3kmsd+A0RR8BmGXEO+qtn
4iDwrZSf8CzlrKYzUjcHePlEU3Lz5rGXYisoR5c519u31y4ns8rYSinQNPPbFGic
8Ky+jU3YoDiVISZLjspq/6G1CojYXVWHMCs4slUJRe5gpl1I2aBElN7LMQAeE3PD
mQF8IfYY/dvQXKV1hSQs68sqYE/ckLq9OpTTH/p8BKQPXwJ8B9G6Y7+ZvgBeSv1N
p2GPUqPJmBsJZK5y9OEpby8Izp51saRikhcJYhmYXtK7jlphqWO+r7mowpQ4GQzP
yeIqx2cWx6/NH84BMEcZaCphBlOtpC+qHnGyvxzKBlR289x1kN+F4VfSrI2HMp8e
ti/U2rIeYOlQSU+AfzUTWqWQxvpAF36tIVWf+dTcOOZ4Njd5JSAxTcVNu0yUijRX
Urj8iboXhBBPKy7ZiONU2rJToEFcCXM4x/clCjtoiejM4vnJp3+dyq+nIx7SZ4ku
7CchdwMQBT26RdZ83+JsSFjreyQ0mhbTZ0fm+RrN8FBeR69eAAfyJzXOyuxWDRrR
gpxi/VwwYKhOVNbEnb5NdeMLzcHvWYkUNUakqk+QoDP3MCvSbbC6sgshgKxvr6z3
jNdg4l/vGPj/COSqW6KqWzMosUmpK8p/lDUCZSI3vI+hYOzIbxnqsfurDy26PF0D
zGKK58IRrbeGhyNFRqUfmSFtnOKkizOs8jGg5hzjvRJaDz/B4wIwCHXcfV/gYtkf
lQCXrq7E/zZko2PzzB4bT4CvolvdTlsQxj8wtS7F80Ko6dH8m9svbsSo92O3d8Dl
+OKKZ5zEVN8uQHHmWlu0UOK1/27dEseVt4BsvXAYBc1sapqiv5AF4YIC1ra9VXiE
BbbXuq6TxBSTBTqA+4uKfFRJ518B0DpMYbOqkUkcM+0YA5W8eIosOGXkgO6arOAQ
/B86ZzR/pYuuvY8OVjQTR84R/bLVJmDVVas3Sbcu8W0fnAhtyIvkeG97JDEbb0Os
pyk+Kh4MdHEFKk9NZd0crXqmC485m0T/BPL6wPJITss+UcBJ2LyOQJYZCQJ72vyT
FRFm3LOWfGEWhlyCM2kT4BpprwtArqemqBaXKwm1onT65sYxkRRSSenlzDcg2F04
H+GFG+5v9LxJBSxINkfycV+/0b5hlynOCylS9czAkKaQel7npuTSbldP4N37svhL
BfzLrk0mWKPFrdX6psDtbigv+YCgow/O0oiHFyoo7s1T0M6tf0bJ6AC8fn+nii10
BcRtpaIfJgsPf7ZCPfvOg7MAy7xYlFn0vVirTVEunP6zw/QGu2kJr/YcVG0A4dYk
7Ju2pbb/GRKXRlLypUMPB9Ri0UD4Nya8vgEIm4SZ1g+QGT2lAWRYs4GtNRUVq9U8
B5xnXXIr5NDatyu3xtWLTjiyXuSkw0+6C8fK0r+sBiIjibBb7lfgsWNZQnq75tZ8
VcgABA8PYVpiGJjVYUWppx5MOKw+LP/91uKmR0Ha9j9DpMzfEwVa4JU6UlkxGU+I
P50W3fpxHoGQbWwIXOeYvcmtFxb5wbBfYuYKIOcRBXWDEDV81Wd5sZI0t5ytYitT
1bR3u/77IAOp8w1vWgAqd76etYfVQuTjpyJfwzd2vmGnIvHomaAoPdahjfSHGdoq
+Le9J4+Lu5CqTKSTTjGVyb5EPCybNYY7v8rQTPsjYXIzcWsfsO5+dLlOEKktASNG
cXxG/xjddyU5LVu4eCqQfPzCh95AogICl0i51vOFDJ1E0B73YYp6VTIjzgOs6Vxo
95XzKm1FcC4yGnRo3JIRW6COSbcEeoB1nNrb2Wc6GSoNzNXfrh3RTlRj9yVSx8K8
2flfHx5ydVADffKc1RzF41pD3bMN+oRDSEys9kZD+yoDMwrErDm0UnkoXTcn66MU
suwKJVadsLdhKBi4yInQuQzgnI28yfpnKuoMh0/fiDHoqd4inqNM7t1x6ECANF6s
LgC/P/QOcENhpTE1BBTA5ySmgMShgERBTJhOW8AXf60tKlV+IYbh1Vw7Bpy7L+HY
w30zTwlzijOOJKkjeRxELbS0WJgLmPAYGTzKVUgUjhFBZPpBDhIYjToMp2/rotXx
wtXPC3edRr2gdrNRUcrfOSvzhCqnHvJUN1oXS4zZMn0gRftzmlFVBVv7xCfExjuB
rlNnI/XWkBcpTa5XNUtlyZE1OmvczO48Y4yhMgpH03k1WbADaRo0XhUB4XIf1cCI
JLf9rwAzOnc/fjelzF3Db+SFV8rS5kzdAcqbqn2HV7ncoPSrjn2iNuH2tjkApSU4
jJTJ4HsPgIULBIwJpBB7MOwWaOUD/TP8RT2YPGkimI+j58fGa5pcddugwtKPwr4i
raiYjKPR1v66BUwQAWXiVNzDJZ+3Ic0DBgMuRRxeHMQ5Vj7eOXwGLNEB13Adm6gs
scBkD823xEoB+2vNVyqr3JRJZWhQFSIS6uQOAKjC/FlIeYFRobWIcNU6FRCIQNWu
0w8gCfIVtRmw5IbmzPwgYXg5jwjYBti70UMof0GTiNern1I11axFKAYXzR2a7gNo
3RM32tpysBpqEPtjN2Blila6f1KJi6zpvgGazUk5g5phOb6H9dYDjNCU+IS/bd6B
QiR02cXiobK+KDi5sfbP3w2NAmiQAC8cDCzVVUW38UO2hTJZZUQPRAtePRVH3Cd3
LwKBAHRBnRazCXvKgbmrV8Wz+vETp/MnuWfvMQ/V5OpyZEMwj7xxlJvgjEfD8vmB
vVrONXw4aCnh1F40BExvfk/X00JrTNiJuz2djLfkUdwemZbMxCftv8f6UkqRSEbC
v1Thc4PxTbdz2ERaT/q6oMMqoHKsS2JaSQCw/KLWce3tUeJHyqQqv+zlYgOzcgq1
Zut0SqOPvVXWAOOS0a7UKC/3rv5LYDwdAyXxAmmZBqV6ymToGUWePpBnqWaJnWXb
cFBNc2EsZfOPfps1rajwOBO5vqrwfQdk2y6Dnpz23KMGZdAHW9236iJ68qu4+mWZ
HeTPecpPTe06cXBg/zaMoDfJO0WL5IPuKrxkfjHBu56UVTppDZYtNYRMxkLtnVTl
iPapdpnX6zMB3KwO01OhwFxxBYQ7cRO0oP2BZmGNlV73fdYslOc9muAfWs8fjQWN
YOyF342pRoxn0N+fj2ipiLF6+j6KirWbNyhAos7O+fDCi9umNTGUSvUXI6GGwNav
AC3+hIAvqukTirL4JG8tJpFv5I1tR6DkmGilvjRrItxGzyTKB5c4U0OuOloQOFJx
`pragma protect end_protected
