// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CYe5euSEeoAdmaXtJNBQjkCsy8QbhtzqGyuYBw0cZul7bUZ4EgTb6S4AO890q/eH
PeugP6VijqG1KEiWZQMiAxjvQwC5L/+2ZmRLV+4jsXftKWuvinmQCw8wNEEoz7mC
VWEwnG6wTuB9qXwj99IFOQ/eFZRMFMfuDrmWC/BKmjY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8400)
mBlE9QCrDDzBTreENMZ5RWTov0eB8oa9Szo0fSvHJfecMalvLRJe2ZGFJMwrluvS
RVTn6e2Ukl2gv7l372my2kVFc821JAtI6PHqKdvJ4sKeMWYcsdq5KWWk2RIfuKxI
u+oI9s5QlBi72vQw9BAg0ZtlptD5kpQHdM1MF31zU7lZvwoI2z85LlYoV+QWuCb7
vL0socAE1qXNi6vnQ+dZPXK7vHhiON07eYKp+iEdwSROrWM9oeq9jSbAyfp/OmpT
Yi1e1VGVxu3BtA7a1tXKj5J8EQgIUlNu/AXAooPnDloAYJL8flHVT0Oo3gU+hiOv
dvEXV7ItJPIZoSy1XNoQJICdXP1tch8wwaFs1g+Qo4fJoof39qjMXgCJfd3xgin4
bOrUFiTeLpw/aWIylJVJ5BfLaiTf5eqt1nJm4Xp1Jg96LlamYuj0natQWnE+Hkfj
reCLBYFdh9R0oDaeutxjB85tI8z7zXX42VTh1yKqHo9W+IFKZoT/DpfdfTG4YR+3
PG34iRP8Y/sB0W2JfUaPmUdY3YqTPSxutY6Lmtv+hxPFh/AV18t5pvACN19jjqLn
OzT1C2DVIbSuR64pm6vLuXLH5QAnE1le8OIrwGYNxUF0gxlsjG2gDoxchjYwdJ0B
HoFAabCdn2Ee3fkqI4SecejZGJbA1n0ZplFzDgjB4pUnPG1AqfS7UNMkh+DbQnEV
mUfxT+XR5+0QoUMMMCeBZnPxwJ7RGcDUa0KFs92rG43THPIb7W5SFsxNQVoYURZ+
GLg7jmvO1TLgwU5gkWrEB4ubaP0xo9YlRddUplLCnsYlq0l8g0BYJB7uCYYtEDXV
qXGQd/elFOEtLrDQ3kA3M4UcnIZU32vAGF2dQQBiyVi94On4hsIBAJxuc/wdt2vs
cQqRHoNAT+84+jnAufDOtQx+IagCRKiROb94YbDe8qE7kXNYG1M/VNkUDJEzqtKM
wx9MGvXaRlEEm7opzayA99D8uG7V/eNmhF0f+J6h0zNHAlFCJWD/d41i1Vpy3hjF
OLYkTihsf6Kdugv26qIEMYb4oBYS3jt3f0YkcYgLE1k/U5dsmFXmmfo+QZe3LsGX
4/LMbbm3QwE03yu+IljPBlGtiNQ/K03gw5eFxYNOtUTkD8u7ghjccB9M8ZJfG+eY
sm7obzCOK/bbio99j/hm+stdVNI8rJ9o1i9KSPxAtw64tlatLg6I38QFihSmSqPS
s6ZPc6UDPqb78G5bYizL0fY02NAQj0nEfVp6sR/Z9hOLM/G1bL7fURKWPLZCb+8S
yN/og0uahEZ1uQhcK0tl+3yxI4AJxzWqkCSsdjjovYU/B0VXZI85RCgj4ekebpqB
Uro7J5UPF6A0lNfCftIVFZkBZdPy8wKssgOxD4H2m6r5wD5cTSNDaXldhSF4xmsU
lYpFBxb252UNWPJTI5l2WQd6Z/2AqtGLriNNJFCzO36olqeH5Xc6FWxBhbxzE5L/
bDt9vzgiKIonFv+WybqQMF0ZRfwbSEYqzAv3Bj8fHUiLz81jgyVC4C27F83t3poI
AUAXm8lAU6sEL/9g0BrDaoXw2WKPIGmkYhE33YKv8ktw9bCVIgdvMLgAQdHwnjlB
p0OiRdVY6qX3WfGQz3LrEL17LvNqCr9DSZl0EV5SFONqrsJAigYBtcWK9WqWyFD9
vylI+1x1gaKR/+IExFbumjfwFlyx4NMM6+8eAwcnts6H8F1/i3RZiRfxmhsv6ZRV
E+2sYJ80pc4xwNYbZnv3ogONy/tKyj2MRLpwq3jM2wJ+6QYdhH667tVdSy51mMc+
elHOX3pFOlCnDXId4151JcZxaXs9NGM4Tnkx2VXn+0Zf12tEObkmPVOYCB3a0NJP
XnXVnrsKghHjilLZY6mmay+++WCJ6A513QiSpM1WY5800FfACFU3PTVK6DCNvoMb
oNGgKHB+zXB46WUC1czArTDICDkULxKOZnofyKrXvuB+zgdi+HeCPQLsf2FzGNOA
VC3Wqep18WiP0olNIsSHTmOorKMkwR0FTAHCCg8OOIy0btphZOOxDfHwoJoaM870
EGp0oBVJ+HZzthXJvfBdH4T2C5R7plsIcvXKRSET0yZwKFECkdE0NxEqvqwJpq4z
I+VvFewyttuvJfW6piu6huJzUWIzQ3M8w75lJajrfWDkqF//oAVvgPEflSTVFWfn
pfnUS7eQvuQVjNsVyUZVGENkzSBGMPO44slKLM3aziVfKHR+RobG3hzwFpBq46NB
2W1+MGqbvT5dhgohvz0TSe2NHK+keyKN6rZztOI0eSUinbCLcpaG4BiRYy3di33q
LKZ2P1ehaHMsOEd4wrufR8ByVYZ9FowQ/xeC0TR/Hc+rMouWcbI65tqIAN+OmuB1
U6gERtUqK5+0ikHxJgTrWN93XPxYqKIs8Rz/pUEd914sSMp/NRpYiW9UKp5Npjp/
3iopwx5pF0bgk8LGH+ODkj5KxFgG1aDDPAQ+3tgMBUcmj9QMHYgrQkvolUEPgXZa
UnIQ173vsColFPJTy681hLKVdxxpVlYTeQvbr7hUQ+Mn7aM2Qf/i9npu7h+SG/oO
S1hhzSmucH+1qc5bjFHxes715ubU/JFl3dNXmuSrAzaOI7PTG7FtlFLG9PsFTBCT
jL7xhs8xxIoAVvPx86PXps00CtTJppmCaqCrvRgvURlhs2O2ssedKckERA/TSPwa
+FFAkfydBGd1i5Mnk9eYUMWCxzAE7MMpgIXdf2rBrxot3F2wNsYiWT44DgsuUTDz
7fmKImGjqcFkvMONb+vEwVbpovCpzaUGd/ewyyvcv3Uj2/DXt2dC5hTLX5m0HwXL
YdR1Jl+TP/y2kxOVcHzmATY5EcuL6aLTklkgW5nOev1wjEBQ1DAOOZM9UXmJG/wv
ZaaOD4RnQao6iR75r+pM2Kpi4nqWfe7OVA/4aP43FItMsIn9i2ljBdnJzcHWSZJG
s5yDJK9uHB44DSYgxcglL54CRqDdgsZ8gOUGrxzMWohOuJtgfTmfV/3I0sL/maAR
FYxdo5tHMlAhfqjw9y7HGtoHFZWIoFhK13KiLP6nPOrZe3Vs5hfvX7DMYwSx+Oe8
nNplKQp1mF8ecWDxMfLiI6eJJ8j8vgmn8wmORZgZA3zlgTMy9YH4P6Npo5RAaoeq
RXJBlWAJ9qigO/DRWubcIGwU0wdYkr2wDBV9p033Sul0DnR9hjXZBAevr7YNh3wD
sBueq3ikH4me4am2mxFrY7ZuIry9Klp3/pcRe92w4V/WJpVoVjurJjojS/MZKEyr
qIRE9vCuK9VKm3dswCJJ76Cws7HCmfZDQj084rPqCFz4eAMuJlfghfQODX16NAWI
p66MUwFVgYOptq6+5W2DkFSSXVFnGn/Dj6saCnDl6bLCW6H+lxoN1IIw153rOCr1
TBoeiMyewdeTp4jht9iAq9u080v1krJiHi86DotS74WZ2R3lOxQRrPCvMKrIi8JL
BE3RjhSaf4jaLKhCztE0DRe9HN2tP2amcDxuYxXRuFh4Ld97vMtOZzZ+ae7XAimF
Z7dm4uSQcUDAhCnAE2YtDC+PTXIEnQkkEX8GQc1+7gomv6UAKEdmYqe7oPhE4cM3
9tNpOVX5om+N4o3HSUvwZ18DCw/MaXez1LbY3Tg2tunVdMADZdNxp30522WWEYw9
sa/+908I17TQgicj0h3nfRbFhtfijLztfNeiNAXx6JKkIozRz3sJ/K+IDIt/JPrg
9KUtwJgxRaY9omRgtD/sk5AJ2G9+xYo2mQgJLMwekzefDdDUiYLQkwmVObR/7Ssx
i2RdxkYQs/xWPfIsCmFlXcvROMn3iWOXdVahMnm/5qHW6OENWcEVXTJvgNIZDfUW
gGEvRcJUMhu6rUUQuuJlcAgRqHdkIQlEpAiHMP4pu2ZjWVFH5C2XT/Nlq7JzjdQF
GsDU+rX4xKRzs5Cex27qwyjlsWBywCkppQEkPF9Z8RuwU+OT+jDpzpZ7JdtEF35Z
dQU9OJzpc+2kT79V32ZHg+rV2nek+RxzSS6/na0bk3qedk3gkgR2bBwE4+XMEsns
0eUNIYPsdtpr5Jr8IFEYDgBh3gMsagVwhlWhJL7hPJkLRNDZTBykNWW6OW1GCE+p
CEkTMyJcCZANabrgh8tabhUEICiKcpkKC8Il2hAWU2a4KIJnAiCi3AMnh8QHc8Sp
NTsDqoFKJhdinUTwCvaVD7NUDd1Iywt0iXv7M4iryu9LQR5cTrOliQmSzrxobhfw
inYj6g9uuuSVnlsqclfxenVXAOFSWtitz4wVEyJL+BTIS1rshRIjlfmOi7771P7G
vlN05jy3FnbkAdmM4s0ryUWsRGvK+TMiY3XixxCqC1hIcASCd4kVOzQbGJIV/F23
7taA2CgzzZaGB5X3U7VY2LctWfjbC1ebwK38k0k/JZFighPUBpnzH2bT9bJ7AZ9s
u3cH2FXMr7CB0nUbxbfq1IcjY7XqwAxGLCfbRxKpeqwxQCU5xHGTdVm5/YHTGSHn
ZcYWSU6HNXA5LXUjHBAvbI6cGCsaugmRvKrCQHLLREtm6IUcBLngGjUKe2OXbXGn
5aSqDkHT/nXkxvX5mO+xMgr4bYjZ3+dFit9ieoGBhjL/GxZ6PsnIv2hWdNhV/sYI
IucUzuUB3A51j1j7EuI3bABsd8rJSjoZXhgAjdmpG++B7DzAA70x4EGem+k94+6n
t/SAKK8EFusVxdEEmPW6miA5botldPMJvgdbGvWcGAF7NIjs5CdwlTZpQ0VF0XYC
+hFlKtNx12h4jHNmw+qL6t51onS442Eu+RIYxwCEc7HriOAUKscAdcEq4obt/tFR
jAZrQ1vvz9MRSPhzle7agRSok1qp4emZ/Ymh4da1VnEACjoYlVG1jy6OLqWDlCLj
Qz+DVzWdZwzOhFXG2uG8UI9Dqx56cg98T0jBlodQFkSPjvlLeiYCgBNFUyzlnwJs
5o7l5Xnsfg1DO806PRziJD3HNRWZbBc4aG67ehKxF5LGqyVDaUN5ZlEKqh5d9u5N
8ky6vh3c9GTxUomGo+qApJ63d7AvBReXkT0UqYthv0CR+D/VWEhxp3n0GXIwxhbV
N/8qeW+d8xQaAFo4+cOF9nH5KixBhUARGeue8X59JM1+HTlWGA8NZaq/MQJSJAr2
7HKoCo7WrQS8umxaQCWQ1wJTiXRu/GkU5aiYwhJPbfXMoAFrkWYjz8H/mB39HA+4
mtwbfXXzpI5qA8COp6XldSC/+U4LAJZAEHDimgEVJnMR92WS0s9T9Kx9QPAq6RCj
lJCL+HxK+rblQmpjuqiyaOJynAS8gxynPSjxRJDxn80fcE/xDfqmt/CIrRe3RF/P
S9G6Ojm2Lya+aLZiK+KfUK0qgDJbYmh3IkouCD0BeJd8wvBsDULLL3cbyESf9tvP
vpVKSXIuh/mUud9qmkmS3ih02GPHRIcusVKT45YqZL8T6QBNhlcrwhJ3brTUDO+h
pmnzHKMuNBE55Rrx1hQqj05VYhwZ1sFDrDochpUa6INMd6K/405mHJ2vHqc9I47I
S4jcp9AmrnnMX1YYnFdTwNjUdVD89UYTcZvnhfE6DxP3ZbEhwJEggrJCgeaodtEX
t/pA3wzQ1wQOs0AhXjxXm8h/oqUUB4SxztR8bvSsCl8GdXc3PA+okR/ftjOK7Aa7
kFSepPDQKTild6jBcIFCaQOygWVXfJm2+Rh1J0LnMS5FKvoYzYE40TlilHNOwsjx
QYDIq0NyaJ4x2NBcrS1A8gvt2MgKI5yYvZRTqf7qYhH1xCy4M6zr35nlt4Fyt1PM
NO3G6o2u3HpG0E4iR8m2n/vqZ/AgyvUGL8Eq5AZJW5JwzKWn9ya4xbbY0mU6jHiV
oPb1gt02JgcDuQ9OeKT1GxlEXQ6ZnS1HQXhvrdNFAa7plzc5Cba6rzTeOaA5odeI
DECDUxKubMJSZ17In9nRbhvSCDdQKk5Nw8NmGRrAaoiX0U/D/jE+n8chKHbcn2GC
1pmhQLmWEMGCUbStYteLLyxoD0NTpF56d2dnjxrWJF35wJ+pkRcyPRmof/xPVrtw
HUgctMfsugACzfW5pYy2a9W/EMQRoyjIlj+X8N15nm4hJQoz3qw1EsbyavO49Yh/
AvPL5BWG7wrBwo2LqehZPovmTTk7cd06iUvvl2qsm0C4/8lcSLU61afOpkWUhALD
gkguiLLzWUYMs4buK5v4FvxJKxYQAbi0slOCTb8p1zZQacxS20pJY+OVhNW9apgg
ONBst9HSK/SyK2FXk0TKblY8kxwoVa/ko8vnV8P8c95I+kZICZu18WwwIG6jJpkC
O5Gk4KYukU5faLlH+aUXntqaQBZTwX67RPaGnDjVlqJFT46vHFLSblyve83mPhiT
oYDQ5Iu/UZ20wHF3LSfsoh4HEtSP+nfdLnLPrt2iTfRSJ0ZP33I+l7V5ucezrkVn
SSTkTtK4e10l+XZ0fZirqXi6p0VqFYv8AB/Ha9L2rVDwW6FROshiUvB/uSldAb+O
q05QaoAINLsjtUah1CtySMeImlNp31qQMUPCcB48ToUkrr4IkTctfUvw8a78eEVq
oehfC7ch4WMrk9N2dPcLwrBuinXWas76hqOBLAQUWuBU55niW1zuxmD+N5q0TKUH
8fpK63eTJq9Ox9Uf7gYU/8XRkOwkuNt1KWCROYVkUDYMaoQBG8AC2JBtGoafK62U
h7jajuszyI2FdfnbwzbMDRdvrXmMsjyjZ1TW1tyJHyH1CjKuc1hRA9JJ2zLM4QNH
YxU5yzX31Pi9CZtM6gCE2kkDfFQWCfXXNWF+7CPzXr82EKfGMdlN3ciMgzeIaQTU
F0bkbYS7Il1GvCwfBpUoQy/oPhv9u49avCpPP7jrHPcIAbLvYSYSzvQ4rsbhEY0U
Yh6/Sk/jvxvbaeZbzRw8gxgVXfS3ZRnMde0VlfyHZUDNzoXr9dTJcvnXeAazfUbc
mnTU4Vu7XJKCBj2CwHxUMUaxbAd7SkJMYB6G4TqxnJM17JgIFD90QFkWIPylM/6K
yOyRtYA2+TZHRVnT8kv+MdPZHv4Q7umN0nV3Krt4Dt/M7fbUuhWI8LlkzTFLaCDp
ZTuYb3QEbqOdeB1LDE4gcjapY0z4ZXxQ/hBjEsbvkYpgA9uMR2kwaDL5UvsyaVzO
rHf+GM2dHz3V//oXl4J8W2e79owHdKosK1acIcFUVdFGogJMH/PqMMq70ARO52oJ
29jhLScik0vBke/0Be4SkSqoKQiOEGGCkzUo0KEz+Fefy0xB31tV5Dl1m0JhXk/5
OH61Ka+ROtaJ1cqTj69rzk6gLnoYN16lg2PppDBkpq7yGKGMvHIIwu7kdz3NUbyj
ETBVF1ot6j5Ux+oLUBs6Xn/2Gdk+DpYRfaaOh2BayCst9IbBURswmDuq7YRsTXU9
Hogv9fpjpIJKXM7PNBHQqIroq/f9z9CI4MO5hxgFrxwvLwnotTeZXG6yQkvt5doD
B4SoTkKzChTvxbeDenczAi6It17F7uZ58nG2Wv9Xgs4jvsYbNjPSdNSFpjz4+VJN
mjgseXy7Zq2kWOy2KBFmFUG9moPeqt1FtnQL1EqWoyIx91Ar5MFxGjyunqw//BwH
tl4h8I6bilsKZSGdFXLcPK9x/D1iOPpJPeV0wKBMu/qlqPxX7Rgi/Et9yHsdo+W0
Q34A7cGZlX+3Y3gnfMutx+sVHEHEiln70ihskhJ1YolGF4cFUpNX9NnpR6lJRxJ5
Eo5mXJAeZyt1+uKB0jzcdwkelYLgnW8LrFGaU4NrlBb7UgLcXEtNmGIWyXJ0f4Oh
j6q9uuV+PyTkSyvBHYsWUHmwYAkqzRBeMQtybLXqqNyf80E9NSmAiUOmTDybhsSF
2kK4v3E491ummz5SRYHNjSOhringEd4MKEGPSm8h0s3dGD3NqrtiQLZpKCUUQHYa
yOSp1CVauD95A1TC1ssJE+RwSTKo/hJMfG1YKjG7EQC59QFCvFAVmx4fZrf1ye+x
aSVqJW0/bcT1WcDoCkM4Q/BKrZE0qNuh8KxSZmemnReW/ko2u9laDWa5entYcBDk
gEki5NJVUN7DA2U4Rt4ZhxvAEEOYxL38TUKkeLozvlQvenMScFQEkJiPqFydoHp9
icAHXdKGizh9i7hVkrBchBaZV0dZ3h0Bnl23eWlf6AfrjbR3DLPxtyt4pOSXD8DH
OB5T5YF/kbZ1eNXljeEotepOUbN10C2+/iY/9tJI01puRzykzwt80egzc3mR/829
2eumKtN4pvL/mVMGbQ1pvo1LS+pTf/3lRCfyao2w9TxoWN4Lh6IXZvV6wr6aZG4R
pgdP/LMK0JuxwWQ1g0e5urp3we4ZEsyPjpEV9T64t2yJiII6KNkMUvZFaq1abld+
KcsO6k643eg9zB1HQKwNTi2qGLsK1XmVmyofBImVpQ5gqkxNQBhhBmkSG3h6KpbH
fA5g/jjimLimLASKK3mQ4H3t/qV47uDSz7JULhKMDpL3+9LLU7BmGBdzv0+8szBZ
dydZfuge5kycsmW8L8QtpK7oHzecvqxJDHbTYhpJmEJUKfswXF7xuCx4PJFlDqqw
7f6YTGc690ba130BWxwXo7xnOoeOp0Fdzl6+Uli3O0huv+mT3lrAQ2BSOcOQvbn/
gnkBdd/Qdolg+mSeL/ftS3Yk+XH5t8jI3WTiD5cGRqyjI3FRT8dJDyvVfPCLRyt0
MppimuUVYJn+k3qHtAPyEhiOexSARpCPmiyFJ8uA7knNyggfA9R+SysFewxOP89g
kGDCoIs20hRjZLjPiThyuA3H9EoVOB4o+e6yxu8VD+ZFjyi2tmnQkYIhW7yxj0oe
nRYSHh35lJJBcG0JbCnjFTUtc2l4FyFIEu6a7H7MNqVGUJ9IhrdtR4eqTZoILy5X
648g6R18Db57YkUhxkIu41xlYSnvAWuUiKCvvqkL9iWHWkQk/4E8gGIPvCvOiI5P
yEABXZJxos9xSj0HRYACyd2CfWfuNqmFJ7HZP6dlnK/iBm8nbC1snRbUDjiUBZfJ
ASE2wwh9808w3slsCBGe9By+dOxT+//YrKtdzBCKhkwwPteAFipJ90eTTSmQVzJ+
S8ditRdNz2W0hSsef9C73eharUNJToEeqezchuU/XTOXgSTYHfEqnS7nLPUWXnrL
0XY4gvbgtKqvLgoifh/PdAvN6D2mnSHEHe+Q1ABvrx5WECcGl7zLiGg8Q+3Co5YX
s6rtU5CRMNrjIgCUFvQTdjsNsEtKHBc3EaQrZGqLtO6yPpAb9smrh66+gcxux87n
mXkGiiIOtA42uZVzrps7CSlVcegoXxQmTa93nkarSntZKulMvKksslLmIFtBfbKB
+qjLxj0+YR7nipM8bB86adFUVMW9Ioya8BktCRgghiRYn9rF1aCqUW5MYbQEvyPT
VkAQaGT9A3fQ+/QM8oT+1T1ugDCXZP0URSBeJD/OsCEA+X6YiXzZvuAbuvzrFs51
pRiL23tyccL3fFom3GdULba5opSsvjkG41ExlCW2A0CTtadAeq420+TXcMoxLIic
MsHFobMnEQXwMVIK0anD+CUVJDLUu8nfyaE2YF3FF28P+Dyok9GcESfTeSFMWEdq
xrQWfKCz7UuYPrnWGo2g0Mzl5B8qp0a+/tP66fsB0qhzuQp23LT2TO7la+XJO5Q7
ZUqYIsLTWgleeGV7mM89MugP+fug4mSd/aQkRqxm8XfcQRH77O3Dm1tXy+ef70Un
R6SqjQfwrhUE7fOEfwKDxM+6VLSSFZfp6RqM+3lcOqQQtqKmfFxPwJ2CxiaCP4o8
OD9EAc4VM7qreOEFh1ACbKPnfhEF5GYx4jZalycPMNw4UR9RdIDuq/V1sqtsHZuj
pMj7wuUvkUF3tWNl3Fy5g9Vmv9qyURXBVBfTUhTSucHddGn125rJ3Es89wHHEHY3
M33Klzuk7B/jx1D7mxmdb36LcgpGtqmmOLhXFVxfCNIo/POLhc5DQLq0Jr9cAbpF
+XUFabvzl/bHOep6Jj7sPWixCJkIF6hc+MU18wnsyiZzMAehOIEdjJ31ILLtOtdU
DYFOS7eM2k7GMWEdU33lM8j7LxKARGMRjmVF2SImbSAcI/JyMe90Fii7a3qgc9p0
KJ0IZ0aDTtBEknd0fLPuKAzUhUVTW/ezcPjz6k+ABaSEAR8TfNcbrlqAibR1X5xw
Dr93MUc5Tjgo6+3OyTMbU1oF1uVEm7bk00Sdobxj6sno7hFExHSwYxe9AEAymcwt
0IVGV3VI8oRuKJrt+tfgw7tC1/8UHeR2TOOhxJT3TXcqPEd7ueAznLNDxvEUhTiG
UD3xXaIBPgzZ8EEIQQyKo3L6O36CSRrgivpSPR6CCOhi0I84O2hdXJcdAkR6TU2A
slE+F9J8w4YWcgZfWTkc9r1qK0/uaABj0SGQOeL2Km0vt59g0yhW35uXElabBJ34
3S1EkD+GuZihcJY7pwJYQXhkHuGsthiuUG/dfcTfR0x0rKC2qorcbcg3u5yJasJa
tIqaJ4O2D8BQi2fLEOQuIdHOsydJ2afiQZYQky18cczKKEE+zguXuJVPN2u8kYGv
5Nj7uyVe5r2o7ip1AlGpCn1nIbj9Xb7ubVD8H1kxOAcYd3i3CHcvX1uonee+5oz/
mi67xpmKLyVk9fk8j3n/fEJjDN0te2eeTzMFwPHhyOCgrxH+ibPItT7o0DwsNzyc
+NYxNz7rfrsf7a7aI79evZ2En5iYlxkact3/7T3lQxOZoR0AtuOUaJFy3j6okPeY
PCrdbVCWxZcazr3LA26kGFWKYIbF5V/0kdK0TvUJq3tRSxoLHw6FUi/83NnK0pj7
NdLWLANo7D4Cw9JzCNtvD9obW+vKGnL9kgFozUC87X61kx1l+U9ztB1WJz1r/lwo
g2gCx80BQy9eLyDRvsp7dSy0Cn6ZjzFC4g4/+X5dZlRAACFSufTVrnW/ZK2hzWKW
V9g8yWJEUp3/DsvJqGOqtCNZebbtCZlUymNES6c4IYj0yk314LcM1Xlef22rEe+P
1w0H9PviUZFV2zAmnmDpto/IP82KSuRO6CNW8tUL3NBn+qoIP3kVqOBQnb0LxfnU
HbwfV9bV6rDTWSRytqiYJed7Fe5gL8hvON0X0SvDr0f56BOXW7lexEaZyZEAjhG9
dcDoVd8RxW65mznyC969ifNsHebTjJU/eDobTi2dG96DkkgJwVxRtmkHyGUNeyVv
pWCESzq/E6/MaTUWdQNxUu/6as3fB2N9FyQ2YUUlsuVEIFnHrQjHKGtS1C2CX2Dp
`pragma protect end_protected
