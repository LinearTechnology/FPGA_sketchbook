// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KR4EhdjZ4V3XmIlakKI4cE4BOHmfS0imAwSpAAmPfbIQORimaI/K97tqDHFcTExp
tH+Fi+VtfKtU4+U/FO+Cwo+LEQnkmxcvkwUjNQgapJQxJb+UneHLdQkIcJPAU0qZ
te/UnIKA4/X+Od8tosjp4BNMWudlC/Qa8yK7UHz6juU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12144)
SpDqtEiGi0AaMvhimx6N5tuRfHRycAoZv1pDIs5N4lROr1IDT7U+W2IYc4B534zb
puAm1WdVDHFgwiWeue2rYSHTpQEKl1qXZNCflPQ7DX+2fcpns4EXcCyAZecNnjJQ
hgwaCpiEtCoRJlHMjzthpuyZRcjKhoG6OaFQbhx1kg97ySSYxYyBK6EZ3fSNQsSR
RXWFungcdN+8C/yS2jFhFVEiyZG7hWn+W2RRQA3ZAviv47uBPIgmmyYuZz/2o3vs
RXHdTK2unBcpoDsopM+EqHjxF87Gq4fwU0eXTp3I4D1Zo+XDL6pA0ZsjDfq60B7H
2I5wA0Hp6M+SCqGKtDQa5rB057BDCZhppj3K9MZeiR8TwWTvVkYm1fMF1BLhcs8v
oAK365kRTk1KWo7L6/RoKCXq0SdFLZWbtw+ThD5oMKVScrc0EBubW66dN7oVFG11
7WD7PE/1sEmiIUZ0U2qmCw6S21E6/po07yg9EVRfOU5wlJ8H4G5VUQtOlvam/CYG
cXMeeExF6vPsfqGI8rDLC4xTJZVqEWwuwyzefN91mn2NveYP9ZfgiXVKieGVVZcr
kvfMZ+gm9ifVQU+VpfSVAfz0aLWUKZmxvWaVL1o80aXf7WRWFGfH9sRiGVaQDT0G
bgHTZ9uYAMO8M5KUWgNwXoD4rfsg302qFQlrY2eLx5gYJvUX34I2Tjz545BQBBnd
Q+FuS4ZKcirUOpEheHY9wO6Yr7xb2X43gM88CePKT17p+E0SPaWhWiYg9QruLDeI
AruutM6WymeOun7WL3twec5zgBtP4glSOCgprUIMACly8+UfE6wLplUKnSZRxfyR
cgfJ9e3dvaJ56HO7l7VIMI5ulm2vgxsPHB/tBZdp1Xg6Us5BCHcfX/QN5SNOe3CM
qyqL2jrg9C6Z3ynoyBfUVzx0QrJJrv6LyiLfBZTOpFVtSI9DltKYmWOcuhH7xIdn
tZRcPDRFe2EACXQm8CUwiuYmr9Jq9IKg7EkwRjEte7qqCYtsbe5klDiBs5QpDI0j
aWe2E1h0ej5XQayVvzQOOKufLmHWNAcifJModWu4+l79rSu5Qwjm1ji6h2B+EKMv
6rEptdXZrjtSqAhzI4IhKtsRf3SRe6UugpNRzlvYsRXUW7sIquSK2SOiNXZvUPsm
tsxfGUcM3SsidyXxLh/KpVO1jT4jt2ZnJj+lMupTvROmF2QhrUvMyi2RK1KynTAv
Altltf+wAp4pjujd4xvlhYhIGYKwKGRpLQleNFcPs7vNlC8Bo/l59L0Ll0ms0CFo
qtyp4ygNiP1Qwoqk2otlLgFIgYl5oGSOhJ7IfvZ3mMPLSpMeq6AFvsHc3wEWLUcu
ZVnfDR9fS9jbj/jNaBxP40lZYowklr/etZ5ZHVfudyBexZyb2qrlS9dVJ7FpFzum
wgrvhb0DcPqKYTLetBDlF2QFsxGvAjpzwnBlgRc2s4+6CoEeD4daFMNYWmR9e8aV
iPN4Y6GDsvKdvGmZDQ+/7ix8CxBlUWkRN13kG9bc7duch+aEP+eaOswc9vh/ms86
ss3wEBNbt+EEsDfRY6h7qZocsnBtcfVXfUtsXKmVGL2HFuWL7VXG9GINZF1aCgAV
iVNZu++cGldgk/ILZQMfypXCGATx4AfYSRJVzxPM0Iag6kzPoWOuK+FggH6RLfwz
rchPUYmL/TiYTsJqIRITvIHfAiJSXAcT2ZZo7GkVn/7UUxWfAEL9qwLKK6asPK9E
v8QsgtWNnEuK+GJlw73W93AuRFUA2WH8UnIXUsxUThY6wZzxoiGPFIbNxQeP+eh1
PxX5ZO5NrvdlWa+TNrBaFIBRqFWGTOFl1nvaHAV3KsMV87qqS55iS8ZNHWrasfy3
RhCwnNr+YxiWEQq/WBePFQvuixcr1hiIP2xL+4vW976oHGAUpfJuZuHW6RjixbwW
AneyCUvRByNHr1jXklAKi1yRv+47CI2P5TWxPWLfSGSg2EyamsL45ChkfVflSsLd
ZtfahoX8kbxptKN47tAbL3d3nS134XRXhT5u//JoZ9MODinRE4945JUnhxV5M0Wn
M9lanXuoCZbyDAoYZnw2Hw5G5sq6hatrUF+ASSwRbFXkSqoRsp6sqRtyYF8vo47+
XF15ERe4DXzfgvPg0GBLggTz7tstioe4CZT7dXuHpspQnKEN6ZYXUY29e38ogyUR
78QZTh7rvK12a9lr6lfJJ1G3xQArPhAsbcHZALIsCGQSUVlesnX0Zl7bWRruKpRI
H7xCWT5Y3fQuGfRKSCOMkpPjB4y7FyxYiWm7v1RiUcCQGGrHDUe9FZhItHUHFztV
z33x9n6cPlPuVzPu4OD1rpzytF1uL2HHv6zF6QYSOwXdhB+kiJzJP8JC4fIMPZjc
2MXQWHd67Pznc40H12P0OCgom38sHvWJg9HRYCFO0YbYcyxpSF4sn8s4rLgyn/1/
pmoAoudtS4pGIttflXfM0HqihzBdZmSuWcctgE/yJWRjtynn4//QWKJhE6bs2GTl
aFzOgH6lylJdt7pxfexD5vSd1Y2oWT4IFHmzqf3chORlrA2e6buchoEoMuhfv79t
JUZLMn+1aJxqAY+TFdRA1Y1BO284Q0X5ub/28oBuXyq2lkgGHgWNPqpokLrVL3ql
oOaqUVdEJRPUBr9GBybG/WNTm3jZVaGWSVB3YD0t3vmhTWxUJLRHATV4H0MEd/To
OmnOxrQ0bSUzUyAo5dovELEC2mQeQqWWHbuPorUsL4i3cwUBE6i+8tFNCkDj1ojO
kWHEncbhIQXAFPKkIM05tK4XmUHZk7AdU2DVicz2BYkw1Jtp45eN6l5tAdX7Snxg
PV0y+G4EwvMXNLvRp8o9hGOFsn05orxoZBJWRvK/n9kSDukgjzMb0nO2oc+bcYos
jlv6CA1l6BL1HN7hVKP2oyuJCYyZM368dAQmCYJ0UHUs4oHtDK9s9Fj0skuIO6ds
z10XzVG053PqpZ8cW/lqyHFSyqPgeIN+mvgapIc4T03L8hX+0+j3DTbd1AaGTSxW
WJWJpOoSHAsrWo23L/dKpGGIGg7rQML9nupxg/LXCLzrtAftFlzz3JqMNvzezK3r
9x3zbuavH+ZcjPu752NI72A4hCgCHEKsKtW2SzH9UtI0Uak0fhTxkfYmpAtfBnOK
JLs9VkvJS0+dl+tY/nR4uAff5aiKR0I13xXaeE3MFQJOi8nJqSg5/4l5koZIprFv
6zt1lu83CvmXLIs2CLhS+Fvs34lgdSadZ6wawwMRCgpzpyL2e5yctYflc1+5Or2q
kTKuxNBssVPqQGcQHPzfRNrocX/O3aA1VnzhsYVNN/WVg1WlQnb6SfVdEIpM9o7+
BBytDComYrgDeqal2VnkdESiloy3URsg5hI6XtvqsLcx5hJKpwzcFpjmzmjEJIF+
Qo8CZUKCGnkyLsnXKxkx9iSYEdPQfzHnzcQlTSWcShSHsak+IzhgNEL9nMZXdQSp
NNznU8Jg0aC84RXaPbB5AGYqu1SQD0g3ZZdHHQjCkRueS4fz27+p2LkabU3jHQmm
VWsI20lRfXu074NcaBP1g4vRuc3mzyp6kdlZ2wRiZc9h7lctMTtCMmAjURB+SyII
eqgElQaGCSHF+jcZk+OeE3BtKYaYxxC6fTiANtUQc2RgyV6MNCBud0D1dhQpVJJ8
4wH0KOBjt2JbYH1Cmw8XYl4i5E0NrNNSX6FO8N7R/QJg6zgizaiWudHcxB7t4RdP
5cr7tQOGVTac+DTcmPy7WteIlyUYID6Q0OnJiJdvvYMdVI5kizTtE9V5r5Zr3A+v
5dAYo7K+ARB1fVF9NEpUMeun8tb8j8X18cQZXSoXHnAV1jxXGZu9Zf+nXdM936s4
zRZhb2wIKlXFWSTxoNZvnR+PUjdnpPdjUbwiy3cjPxK77NZUHNoCeVlQ8lVgOq2y
WDKSUyKckJbCWZrGEpBqBnrHLEBYdB7APqoEGefY4DXoQ+kmfLwB7FAfTtOl0fU0
qluMs193b3qdVh+Ec7YbFHfil64TWHXasrywrmZBtKlm+04fRR3Z3Tcd/U6a7kPH
mYw+7elbRAzcb9oN3G5fBryJ7X/gg6fTBKpvy9zkR2ETVYjv3620eYhuFyyVdgeY
NgeLJOF2qDt3OnDH40E6O0DvlAtiL81AofipNXiKSht502bIgFyIWbFH9jiBeb5x
slGgqZ8UNSOYVVIr/28IlydFqFzU3a3xHt4e2wlc/Lv0MPfdaKyOZK5cfYfsQ0uj
w/UgsFcoGDqqNfELtHLQUVPJYk9Bt12klkdifXMH38o5pv3oYV8NHbYDwn+38Njc
UYbmUOaVUqWtbIxrex7KVFMLGobU2grb89EtV8gQHIhn3vo8izwIBo4qOP8O/f6+
QZ5CsVUI+aW+LFE00WH4Dfkn1KoZ9xmgxmGSZzSJ0zfMX+f0LdUt6xAKwnCNOSLS
XncmQIEG/18rASLnzbRm08cvPemJhPVraPEQsEXrtKpVU84V621dTaDqtFKnIvLf
c445vQSOjW8Hhwrg7X4aijswYKSMFPha35J2kgHbJmMT6l2jymY1Gu8ZBFfvArQQ
o1jgpAQb3ROy0odZEaddfvywx5mh5SBi2igfrvHMsVIMlU2DwpyY27+UKb2VDn8G
a9hzDRb5sQ8iSyLOxrHJJQFJ14Kz84k1IbsXzoLWA7ysQ/FMcB1r1w6ASzIxaft7
1qW3QFp/OTn5fZ8gB5b7GQsslXkCZJGnTDApf0gKMjM8RoFAXsr8tk70eAlRcJli
GwMr/P664Y/NV6uWy73YoawJ+lpVq+jW4fOseGzbDRjo423IhhrQF0m9qgCe7HUD
O5FeLqCpdz/DczJPZXvj3B8qNAOQj/2CN44ruDyoGdxqgu41RNUl4nZPHnkEgIeT
xq1HNj3THogWC6j/PCCFN3sFJzRTMQhBdTixoEBSsIJKGszZfTqd9Bn0S2BhXZJB
YGZ6c60Is9pclRfAYACqLcC15Zays12nZSl9eRbom43pBtnpuuMmJSfM7cDpIen7
Pnao0zNK0fsa0RCX6zCGvApDewH0m+81k8unmIniXy3hK20aLZyra0J9aHBWedFP
CVJLMf4szVdE3SyDrLP6jowb3+jhhHUQV7RUniu3oNcK7YNWbwi+eues9NbCV3gQ
dzCx8p7w+2GeMTysrcSS/Wdr200edNh1a4LASctFiFO65PnQEQQaQXibjJdLdKxE
uSasnCgUgX6eJN7M1guSQJE0BNfnT8yjhDuBtdXXJv32d/ItcaLyaQHb/b/3/Nqs
GLPaeZ9easnTAL1t6Yd63c/HOAXJHMwapXWBaE81XOeVAUrPnhWSBcQbS+cIEeSj
hpwN7SkujkhfUh5iSNbxHDvNRqnsxHQZqWrVfvlndX73oAwP52vjIt7Fqbw/FKt0
tY8P7i+CDSFcQycsHgTRsDFn4IXPmS1919LSUmAZbYKbw1teqFyzUEsVhHCRQQci
xk0ZIN63KtAL+LB8WEwEvYkuee31J0TIraoiRPAmW3NAaltTt6KxsD/bt0+ZX/ib
aP5bXW0Cu1hhP5qWaufCmwMnZDV0tGs54cH663+pKoBQpfDTRdx1hpyT/V/omWFq
BeNoHsaBBpcRJYDFlNZgPiYMw5azpBQVzsVY4ra1h9yHlGWL84qL0rYA3oT8EXO+
fIw4WPo2lTjNKSqk8r5cgPIHzHD9nYvOohrmCK9/GYDT6YNGhu7QGKGCRL1Tg5d/
XsMpeJ1C3zFv411STVS1b7w0kh/Fw2w9SCAjOcnYN2nxAwJBs9aziEAqVI4QMPmG
7Wky9tCs7B06zXzZtYONUEabwtAEo1gXRsxQdRNARYKQoBxjgoxrRIUbnJgIVgNJ
77ssQrrMVAm7xIhCVhcnFqUVYxnNBK8ThWKlnlL9eppDS8qImd03wRPjyHFJA0Td
d3W8O3FAlEEEDHSAXa03YXT86wvBAsfW4H1s7QvVHp6AMZjyo+d+78eofLR8cH8E
ktCm54QmkLSt8gxHbPrIKCN3r5RO8H7XR9gTnnpK3ozl7nuUE5UOoIuLNFGAd+1D
HHXwe36AVgLUGwi/Z29gV2Kd4YHr55ZGBK7G+oNtpfMjqBI1t0yN9U2Fy/20Owva
5AU+flj5nKSIVvqITbn7usYjJtvnSNdRCjoinnZ7rJzcRaTDWjCPaa3MQ1FcTH3P
ajMv/0n7yBLONMalIIWbreDKOJ8J/fDYOcpkzksh5KCWNmDaq1llvwEDKF3YXVHm
q7dXQk8JszDGu0tNVNG8PpvyjAAo3yd9olgYo7QNIWQULMR8w4FzZS433w1gbjeV
/R+v+nlnsxIbcnR1xU+QlJboW0sG3GSUObcnQ1YyDAWb8upOyEDwiVUAUD6LyO98
ah476wZjKxpDs/aeluTTfewilNlN+ZDJOU8wvoyCEYpYbFaSmRQZAJMvzQ7fVbZn
uBYLFQtwF56UfnkqZA9aLKhiX54r2vO+Oo7oGbGmzz5g3v4sM6W0KewrgldYmJ81
c5W4FGS0+LcWSRcJ1pcPZlb5/9l9aH8Ps1ZxZ2iBjN+Gspo2WHUBUVGFV8YZfNmW
JRco3eTlAPY6QIypvEvxvE1pdQDPlJS2Fg6AnauIyTJSdfPrePIoEXorZJ+W1Jmy
8M/6mo/MCez335xnwGZ/4zv5blF3JCvJ77nfLjVGJ7MUl21ayrjMGlq057lcIA0j
7WvJtiRGrWR2dzFzl/QYxWnU0F6jQB549YOwzZu7IZj0M5AIJ4CPuT3xz5fBKdT7
WdHvrW8jFkj1/67nhCbaMKEzlYjvKTgkLPtChWscroPYk5H2qgFoFpS/AJoryZGb
utidSB2N55Wt6cmTOxCmEaaWHjDnkdFUVAIcqUO+1jLXyELGrn1xRC/MxgUn2CHc
KfpQaTiMaP018plwR5IcjO1FdYNWxD+eweuBNk3FCPUL8MQovpbwb3phNgMgyl0t
DVw7uh7QaHge7baTUiNbIj922vjn6VL9bWAk3vifgQAXoZdAE9OUKgmOgbzBgVYT
wTmhBTvgdbeXs9L/b0mAGqkVVd8LvDRJYhZ2AtyzdPlR20VxKW0amUdAyrSQ/UHg
uWDJ5o8i6aAYwayMKtB8T2KInIvfoe+cDCFi0EAv0BHcomzCSdtYn/qEyqaxDOzq
z5UaUewJF9qVI93OXrHwbDmpPzWt5/d2zvZ1SbV5XZU78kMkY3xOUL6YY1nvKz8u
MW9hr3Ymsbi2Pha2bZuXoNvrpPIb6YEhz/+NmfNeNyx/5ujBHKCWf7biWWCYBaW/
dxYODVPol5tGapvqkjTZUS449GpRJSbDR2RQrWuh4Oac15/SPxeuiY9LN0avHo0H
uSH0Ozvnl21OOn9+fD09GYggUp6o8F81qFLczTS3wRR2P+R4Oi/8gifbmWfOdYbV
whiFDaqbb1FlS5ug6GDZIcxMFL+l77yHQtgE0+g8/sNEjQ7ooii/SAX8f0sE24Hp
yiTcrJR4GckzUVOP4X9qTO+MHaI1stPUIsMfcBayqW7UpjtVJFnwGpgY9fwavAPC
OzmNhRx2guHe/AA/VPEVKw3LPVkwlE17L3jvWGOjWF1uSaSEHFh28jGZDU8oBeXT
cuihfQ1ECKxk8q2n2w9sy6WkJm2DenLJaXN/vY8MlLaNZxuq2bdUw/OM9Yv6pDZR
AA5loePPtjaziiZMMGg8mz1DVHdCqgiO/XQXQWV/TcjSbl+DPmoNPYFcwTRNJW2b
NbXkFQwsltm3UWX0jwnO0ZQyygPrfUj4pmA2igA5X6hvi7+H08hFv3+YZwfdskpd
K4HbqOWr+nE72zTn+2wJv75SB+KGTxQ9BeYFQjbMQ9v9fuNLVpzuGICX3TUn76oJ
1T/kioy+NUZ2nZU7DbssqAcUTTGaapZEHIf2WqezzCLb3qh1nVzArth6XdkK6avq
k2TJxw4/J2o7AGtOe4Ruq8mTlm0lIS59z0HxR+EknPBL6YHM0QYT599CXN3NmxPb
76+cOZ1HTbX5E+y6IrBGi4UgZB98H9ax8VgwCXqJuv5l5GjByBOaYrcPItjv3lYK
T5lFsL5fjLzUw8wIr3wEcY4c76Flw/TAMt3m8rfQyR2WS5TkDhqEy9v00Lz1ZyjR
i6g7NQjdmsDtl/z3KDhJXpJfik4FMShmo3UaetZ8a0gq2K4/HigK0eb7mp24AFVR
0R89ub7hkLQARUKwOBCoiS/SAfytnGXcibSAtAJsDjeergwanYPGJ6aTIS0ASeIN
gPGzAtox71rd+iJnQgQwJR4URcaPASrRd3K5jFfN4QTr/YCZoCBFwFm4Aj4IeNwO
2Q0185XTLQ1uqJXNV7lV8suGFSQSxv73IaBo63sNWWF07LfQV9BirE/SEKxR7unA
6nyAhSkbC2gIb+aZdSSCvVtuEKsh5YTCqa0m7kn+TFZrg7pZ0VhUzT/h5X8oB2Qg
qMpzMib+tpOhTPzbZ3YEUfXG5cfbFHf7KJOrCIFV0sE98bz6cfNrZtjXTv7M0biZ
G6Ckav1refYVXAmMdK2qYn4mnM1qyiGgmlcFD6sf23UbVpALVfzWHcz+CY4lf5eS
DIZe/OkpW+nGkoYldw68ouWxFYW/7yPro8Q7eps6Kc8Cp8pAhS7wQKl4rcuRb4Gp
D1oMk/E55c/JuwqAioqPmmUwKseudwbOn2pg67Sa/27eM4rZja1PymTEVEUFnH+m
otd68YBvykxLInfhV2GOryNI1SRI/N/JZEvGQ3gP6OiGPtXS/AIVDkqqQwiNAF+8
ri6juAklWTYrfZvL6a/TP5w7Wkf6GYy99PUQWeBulQGtyZ0347mJzqtDyaNOzU5P
7EsfvkycOnSW0C2/6ioBX41czbGuuACSOXK8oA697eevzVSUGjDYBckPz58DmkoF
U/FhsC36ruT9nvbKvGV6H83UVXE/YaHZc4VAxZVdz+OKNX2F67GHh6sLEqjujfOy
HO9FW/B/5vCz/Q3hFSGf8r+zvQzShvIPNfWnbw/q4hMOkpRWssVGYP9jSE+xU3/7
0sIRNzPH8+/CPkAX+HRiSrrfzUUZQ8ZSKvC9fyBOVDHTQ2SxazbqLt+TWH9/VdUc
J12EpSWQpblGlcEnsIfMUVczYLF6TDEo3mL2fug/3AD+GinztE/Ri2gu5HHpHW/x
ZhlQElD3XVynE21Ybh0ogcPebvPreGwWlGvmkIppcv6LM5H4kLjDSbpBAaULDXsx
C9WOeULtUytoQO4kiomkTCaFMYjWCwoROZonwiPnJOK/MjZmzKgTSaCh65LJG0y7
v3ZTJibZ+xq6a3PtMTIINp6xBwuorXRodAb2eCLV1dUj6OIW6Pmb/OcblGbcHBH0
2FVcTg0UaFvtwZVrSsMG+/6V2sJ6f/mOG5JK+8kzGe3CjfsJfqyUzgDG+AK0UK09
oK54NF/HrA4jSfYPrI3LkqGxIBGIh5x2q94i6mFUzuz/hVg5Z/1m7RCt1H/9thoJ
AleCyNSLe1ndWlak7NV2t2dQtGRzs6x/RsE2uA7Ok4yjycWDirK3EakpTzdWyM6A
dVnfne8plr+ibtvH+tCr1BdOyYjRkn7TsNkBeroRmn56pDAFRpgGwDSqBybBb5S+
UBWdOz6koi3CMpG6ldRQLN19eUblLyGshTVh0styD2MZQ9gABaWqxbONYoza60Dq
gFxcXZBnqO7DsQyHQjCzdk8SeKcddULFbfqsdqz7GT3A3AuGyRgViuSbzu84vvZU
DVVbu+REwd80Wfs29sMdMq5qmr14ICTLXZHDac8iJVKrE270thcjFpr4Cn4sGkUV
oHstyjQbpVSpt5R2spe3XnTUcZz73G8tqimaZ0kLCcUqBLeswaHEhoFxYT8HP2lj
ZU91IlZZIdm7+8D3noVpD5epzUbmz/rmFV87yJwUvNO0ZErZmLoVNOV/haVzwrdt
XBJeFT6OYLTYC/h5xVzzvWODXhF8nDN+V3grgSjdG3jQ3W6hcRBNzG7NFcCkQfhM
jq7Wn7C+QSQiGKV59cMOGOD+Wn6BC5bc94aHkwtdv3OdmHXFmdSq19V79x9JULMf
l3++QvXFpQ2x/IKV0h0FkSfFc4w5ZiLhQGcOJQA3L+E7bY9ng8pkazs1NVKWTHzq
HX0bqiG0EjtUDxqIOc6l7t4Omm312IW8Pq7z3uscRNNW2jTPsBEsHUy5un5vUvsF
kDxOnvC7pVWnXkg3TAlL18+hiwjRqgY/aZE5gm5zo4vuMeIVLjc0s+sFsqVc8BkJ
mzU2NrGxiKdOzc4lAKz4WOejIS41R68kCsX9xjP8iUneyozgf02D0ivaOkGjvFYK
nCaL6mV8k1ZMKskLW7rtc3ALUcVjHdXqy48C+1NtY5m6nl93YjrxRN0nscOWE3wm
1yM8aD/WYODEHvNEhww0jXEyOa1Jm+Ll97ITxZK4+/PTdtkMc2FRe0HVXDcH6Nnx
QhrkOwgMbIxIIV9Sfge8p1PWOogujK/KI/APEL9RE18UeMKK+wPwPphgfh9IJ+5Y
kmwGF6q9o9AxEXlVe147xqeH1hD70zeTE8V2ids4fy/wAyuwlJ0QKkygx6PL5Hq7
YGIqmK7/GuEnadXCtLT2s4nIw1Ch6esg4WlsbaKbfy+euWscGH/qYTgFXThKmTsa
dgF5xELzRg2GwHp9nrd7Gn43O5ZgCjLxVtZOgC16jGCEvj5BZPon0jvPNwRKW8dc
CxNluHUfb3wA1AzNsa5v6p2rZwPWUooD9a+KN6tsRxo8GrrB+qITLt10jO7cmcxd
u0yXHXqSZSM3XhG1MT5AEKJKYpU3IA2LNPh+bJB1htz9R9z9nxEy4FQnrd87Yy9A
NTS+B+HHrMSEY5a6xA6Lf3ryBSQ4N3W0FZzafJdutJIyM6IB8WwxqrWnBCpqgOQd
4wpBJbeaPTWf0AdrFbEmg+cTLBz9f3NbR6dkJAGRL/8Vh7lZcDykmt2gptJSo9MU
2K2tq3KCbsGPXSO70/vx/pWjZEU/9AUMceybLebBxUmCY01dAQwI+WgXWo3eSz6l
zRylSTwBrsbu6wcbY0aqotksTXkPGyFqdlpOMggcB+jSBiJSiA+me93BtVtdy91A
e5X9odSQ3Z94HzYJdTSABM44L3JZG4Q1NZOIcjmIgnjF0E35JuNr+cdS1VXBeEXX
aFjfhVLLIxMmX+wDQzFjkIS0di16LY+vze7LIXLI3e3S2ODrzry6Maj5ocyYktKI
MekAs8Czi3vBQ+rxOzNHjLnCBN4sFfsM8jcj92ri9DIBxmODdaOpndE74/emFahn
NvHbW8oV1n5O9Oniy/bIqGjySPEt4vDhngwPSG9RXk/fNsipU0vA5k+zsWwBZ4O3
3Sxbi+O/1rtV4fe163UrCLVu7B3fbd8IqqE81l9v0YfBIo/lQ1WVQgc1m7lCAIJs
AkkwbReLxMan0K+gG0TGDDGLZ4qWgZ09Jk0exLWoWfwW3XU63U0voeFkXXXlSlfk
Ypt9ElguNki2UYT6QrsgJgZkfBmGSLm+rJkQwvvvk6l43dDSaiOtXZwtx+0hrG+n
5uML4CTEfPnQ+a6xZ4zoQx5jGevPpO/ew4Q02sKQWy0LS43oUksgMjE30uR1Cj34
DvNKqE/hQSz4RcrqUTd1g2ahZ1VO0fwPzdCsQpBnQo/EHIFrJMdBexD1hLn2Ykaz
4u42YcWYqCayAco0CNxOFcfUvI0dQVaxfMnWZjMgCcVuB6tTvTKPEQvCogg+HL5W
dX4/YXlNfqwbSOntdF7ToxaBgrUFTeod2RF/jonlBTMDxU9ZeTkOMnRRaqF7rptO
JEYABdxGu1JbxXbr7hZAaavLpgxsDbldvOp+jXQK7a3yTQL2htTGO7/KKeS6O7gj
Az6T2OgNiBKhsBsb5hDbNaSsA6whxP55RH3WLgW/FsFFa7lPjDbENtmshLZpNJ4D
lGF0e+ctAoFYiWRHuo3Tu/RXdlaCslovHa/fl7uDl5RUZmPp+uhLw97bHnEuPQzK
3HJoFsSkpbwxppNuKuHVQuevGo1eAFucCc4qGDbBBvUfymzFZaxxcxBrgQxNCjAq
3YM5egSK0CKfgbPbk9AtrkSgnuRIg5/dTmXDmqXxpSeBDG6u2dsuVziq1zMlzGM7
fwaQ+AvDrdH5NnLosYfpuRi3elGCqSPShi5/8KOmTCk/VdGM6axi/6dgdXgRks7Z
NEl14gT4M8XkeQVy23RMU5tgYip/Bdv1tc6CySdo3IEO4LdlNYYPm2BPZV86uWEJ
vrwpWtm9SaPHjTjVDCoV2p3qfIgQLD1IxDzeOyqjyBIeBlVskZkbv9nfO1nkBQo7
jVnVy03ArJC49GrI2RBDvgYv24JmkaGaRSUMC/nYk8O0zplgtvtGMQgC+K9pAQF0
xhQujW2F8mxevCovriMlPcazELlI1E5YYqoiB8Mh9umoJigLHltGsr3knVy8yFiV
pXNclj4/W85MQIWn57iLLSHodtVwjW0992W2h0HNAbfTmLr7zZ+G/0Dk36HeioIw
J32DouocX7+yUunNpoiDXCx8qIeTbbGkRTJ/WSR+rhOx05B5lrom23MTbYK/6Pf/
QOXqm2x9pVviEGX7i35ZR5ggN4okroI9TtBGcmQ8j8eFwzLj/gc91skGhBRdnpUU
IPInMidT8+QmsUzGZVQdKo2cDcnzObKj0em6UIdcJpogGWScSfqU4X74h4iIbbSZ
nzFLfAMzmtUuDz4guWQBw9vkMRZ2UC/Ta6EiN8ZsdlsXL7yzJQlbG1COx6wzN3IU
5alLdH2lBCxMHpnxILyr/WdEqeqRe8Atu55FY0QvglzryLGsnZ+RD0WUgfICnBr4
j/o/rnEcqfRXadRQySR0Qk+a2dN1ReL/cbAun71ErgfapfG/39xvO3eEcsgOWoKv
TSgAW/1pI1fvWoElVDArkx1eTp164g206VmKYor5lQn4juez+/VJcvfCS04tXiJa
EbdfCJ8CgrIfUeSjotfFfB+55/ougahtUo8ETOOy0aOfLB8daOs7cVLk/+Hktis6
nSZHW+5wLLWKkon90e0teXDrsUOW5ZZKPWugIbKEn3SdKadEuRzjzJONSRlLOVfm
jSmR5+DrBXC48XtdqHGc7Ie61Vl+j5vRQXIgqmFmw85SeAC+3X01vQJD8JnMcEtq
tpf7Ue0Sb2vCU0CCI0mND8Es/iAUTQXUtuOHhjJhaZMWM6ATiOyNSH6Ld5/sjY0X
WcSFiCMEOlEMaSzjkg0NR9I6zz2KgfIy2pWpehwyfga1ug0qiXg2gex8OW1fxH/+
siJx+yVQY+qVvW4zGmFSvUcKscQ2ksQUuLXIiyZvvylcha1vU6mGH7zHhJyeW88q
6VmBwQ29Gn9HgHAnCf22mKP5dLcabFVlOAuDBI9pmjX4JNttcLAeJdc6CpbA+yhD
62hP6UUPZZM4mAY0tiKUpdKMC/6oTqyr9jZttCkyn9jgd8YZGuOFWIxBDdsZQeNJ
M/D4cFp/UJ2YijxyCaO7C0SvRyy8kbVJFLlkXsGmlAFu4hGKHpX/LxogXJ0HWI68
ijtALBGtuYaxIF0C+avugbE1wZGJhx5RmTxgUQc2wCuduSNXMGVirIya3ZPtdHEW
PsHrAFMEeJha4LYtfxt+57FlHIQ408AWGUefaYqYoA2f4HCKob1thhIQ5+8D1Nbk
LM5r/zOoVb4m/yoPmFwouDzOiN8abzQnREtcYaJ+pUIbelhD1BRi1J5FE7e/rRjA
JxZo2oKH9IQzCbSB6vtoF+lcd0cHxmdISUc0mEfTEGEOC82fzk1UdvS14h1W3KGK
74sqwmICdMBz0CkI6jAxL53ScmxibpVGAodsPZWgZndA0DCw0KfWEq8ZlAjnFTiX
vB6Lxy55zzwJisCuiqoojrXte1BHtqges+vTmv6+3wXMtT8mXsc2+oOmNx2+jzQr
BPNUNTkiOb9ORfPQ4CsVnzg7K8glmuPe4FSsDILb4r81FzC/JbzRmX6sHDXUVkxn
HVkGQJnx6sbSyJzKqdzd1AKaAPuM3R8NxJLKm55BkXQKuZe8vESEP2f9+hkJTSvZ
2b20kz7CfmbOBCD4t2jJWA6NjCKNE8mv/nub52M+bR5OeXv2+T0F50mmfx2tmpzx
4XnePCK/YYH8EBmT5TgMZfejk/NWV+FQxTcYa7VKmreJGS1eCqchyjXZV+U3vU0b
ovvLdyDLa7KC1runndKjHXc/vLHmQxCLi7CIMGCImGrU88d+4KuJr6ixtgyazd2J
u4ViRcDaQ+KIk4t6WCqlLm1pKX/c4AGRf4y0DPGpAGFme43MzFTjUf9Z6Y9DnrXw
tBh4MqCaA+d496zR8azCVvD1M2Vf6Pgp2vraQLDeA/Ukj8eDazvhxlMXR2zyoKIP
hzS23DH9KeZSQCzHLCYpDVvr5qMGT+lX1wno7tyc22KAM1DW6BO0x5XUiB6sV5JF
QWH1oFTBbUqg4TcjYWc3FHmhDaACJNZhDOlQlswxRX3UKMErkMt2SSCLLerHawzy
Nk8b6lCwvqZO2H5wtWiPKjnzh9zosW2KC9wIRgPrF5LBVeGUUfSPaOkoAjZ/gj1K
zJ28/EWQh98PPVp0rG5uncHmelhcZhy37ArBhVXOaYbbSfG8QqlzFinWKkDMiK4J
Ff3MJNG3pUTU+xzajtMocwKpAlc2ajNqeDSeZqqX1vUVU1pM7kXRBrbVBBvbK9mu
n9UXenqMv26V8C2fqds8bqmf1fT3tvaaZ1eWbM0rJjJ2a3Y4uY82OKSLQW6Hxo98
WpKQUg8tj0060KHWhyBoKNxCj3psMcd6+b9A10ab6KZc/qQTPikr2cf0p758JWXf
FgGdP0f3nHtRAc2YoiPlV42wH8SssIGpmJvl9neJIjbxI1Z84EGQfNliICYdOC+p
Yd0Mt3X3Ei44jW1Ct/ovTeVplGegC9yE8Bv775nwh7nCErQtJJ4rtxGaxjTF/Pgu
ysNdZxS59D7gKFgrR0uSYKwk/d8B7xKDWcekQNH/V0bkgBxZcHRbTE2VYT4si1xU
X12USn/AOOU4/HNAjjDZv2Fn4rAJGrhVhmIV0tvZJBu/ELyUUJ7KVBasAtAwOap9
ptl1P7AKu4m8n5lHjqFHV22p6ULOEfwNv9cO/lXl+0J/IUiApvTY8fAPOKoc735u
1Svs9thXOdO3X4HDyo9yyaiEkXM7kblNvEkNemRjjgmRcyzP7fIa9neFe3wdJ0sV
TrZKbIqYvvJB10UiTLbDm7UnJeLpoAIIYpMf6JFbBq+uws6Xv8EOsRik7KmtZOgp
SAZZDAFxrTfCAoDGtjG+KRuGGpg9SHyNrBs5UndjZ5vKdePBlmyyLhCfuaKS8ECz
9JwdoZJNscmDiy7Id4MVV8z/+RDTHI+SgjFBBEIAZDKHn917cInNQFQSURsh3F61
w0pQ6Lj3yw4kCVax78XcIC5Yz6g6+J5iZ9fWcFX6H8Yz526TL6x29mF/B3wPDJd+
6d3Z87KTKBgW1eTDFY1mdEKkp7facVr247oFDl9IxHhjVktEZGMG5/ENjUMQovlh
bfFOEOhttdKJb0EDoabNiCgGDHhNmJYIKSuOErSubBc0IkD7mMvXpekB1UPLtASY
RoXak3wPqvj3oKy9VXUs5q/ofrUUgqDSirS9XZR4qdrj/oSVlUNcuqWgywXKCPNQ
l/UNE5NwT+hWGVo9hVqHnd1XmXkyAoK1ZDxqFpYZcHv7IwTpH5lOkiGLC9EoF1FJ
XUoynV6Hd+2Gwao5uu2TWLPSF17epLn8LuDp0yru3WMagRWQNPlJiLnVsM+4uY1H
qJ3c48NiHV5PqICG8wGwOEMRqyBuCbegNZhZpVbl/gM8u3ZXTZYWmfP+iKbdAW2o
SNh7w6bknMc0FYcoZKqTCniSIToGvo+U/CAs/j1M02JuUShUuvvu4c5bVGQ6jv8X
8FIK/KxQTnl1Yl0u2vHwD507qeQsyNtTEUuNXMviMaSDecPK8huL5lZjtf9Aczcq
1TuQ0pvbPY34dFwM4bzpaatQXShxWjRRvob3vDhod0MDqA4ZrXCY9DK1/uh7Dgmn
MDcv7lt3yLFrt1QtcdBlGj55mzQkFqAUlhtveDVhnSUY4Wx5jY/QhE+oMXaAzYsL
zfTzbBuRp64HbRfWqQGzz+yxNsGj9C2epKZ5BHRINfQGxQFVhacZ+Rra2yh2uZHn
D8PvRUUl+ZnaqYuDh7cFPofDX6ts/Fs2WvKShWuYEnICdr1vBNLPWv0vPEoFBsYo
Z7GjE4bs9stC10rv7jfSKgXJS1ZDLoLbuasqrDZ0ONWXK/rePPwhdiVJOuKeiDKr
`pragma protect end_protected
