// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qKh4D2C2G6POT4V4h7fEGlZ7QYNApAdLxp1ck34bpgqzEpQkpKBr7791o2mW1xfF
o698O4sziphosRQVPL3+oaO+cEChJNo2+hfQzUbW2A3IBQD7SDSshhHx6aENgv8u
RuOgeQYanS0W9F66TsBuC7sCqbiNkGBm8PWcPsrwx5w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13232)
NC5Ku6ds/NyD8/HJjeSFgIxcjS4BQeOzYMunRB73fw76P23o6mQaZxSWxgNKJYcE
OPiiLxMcAtz4YWiBGxiOvLfg4AHpOs6H+Bkz8T6AxIKBxg7S0gMb91MBlsA+N6wp
t3Zp7cAODfRYTg1HSsKMFx7u3cwfSTgsBTWHqg9S7HNBMatax1lLe11bF7ZfyNPJ
D4qLN+2Io/maLhtxdz1iXPsIFcFpZInOBL8RqokXQKXE9zByfWw+Q1yEWtAD6d0z
b3jg57IMjd3marvwMOjVKawRQ8q7dT1MkQliIzk1Evt36jsqRzsd1eOHDZONVRDj
MqdKzbVe76WPp4pOwgJI/GlaixVl0JOKxIhalnztd4pKsYWzr02mjJBnokKay1rE
ArWGI9h3FhTM7lJ1xvrfs3GXF2h4pMp+DTox6KssHUAzctLBV4EQ4JdS9zS+q0DK
M/z3eOY541uY7E78ZFsX1zxEV27N8HawW8+rUzfwj/ZPuQ528vuKMuHNm1lWCA8p
f/kNF+XFRBC+J+ek9Jvjjo57toT2SE7iFfi4Tgjxl9movUKDWMnts/F+azqQU0wr
g8Qoy+Ej82S6a5l/0rmu0zuA2yzH8ceMEJhx7V8CYDy+vOM07D04UX08KPYPLpDB
J6KTefcOLm8nqZeahmFwXBNBvZO+HeEPWco4DuPn+s+L7+kSy0bIQgJRpkBakcC0
ILaLXCkvpj0mXtZAhd6YN+hgCqxmE9OlxwGye4vkJXt3N+6Z3LL2JEntn0xRW5Or
MoOdBRcfGIrdYYK1PVH/weKJewwbEZHvyoSXufYTDpd28zhxhit4Gqmv+aqo5VuH
+5lKGDKtRWs2altKIcZpX6yvh6OdFKWQTnNBkbFhaSAPFBfIQdM9mnF+Sk7LZb+c
bJjhx0ZTVuURgunFYiiplDuaJFCN2BaHSJ20HwgQoCH6s/iwyJhdn81uArkcWEM2
g425cRMyuxgqJQy2gFTNit28E7LyhD4tCVGVQOrB5t/zTBTUD9Np1c/9CUlIUySP
qnwWSgsxUeX+D+bWGR9OgP7Bm3YEJiq8mPL6bW9rrMf8OcuORtdkFYPx49gRASZ9
yHvYE262wLTgMqcjFvM4wLeKb5phoGfRBA9jYF5lZ1yiqyYKVBJzlESfrKvjXvXg
1dI6YBbv1tbW06QDbBi32CRpz3j+/MBZdQCUozq+/hGfv+/kFenuiTGIQqEXFa4K
8plObYW2Zp1YCwewVUtpojU5++9HFeUeR8DUS68+JyUa/MSINPMnnzJHkhOwoIy0
LQzB6zp/HrfpFqyCDxq6pXPKBbHU9qZYQE6d/GDPd+LZkBap6tBKg+A+PRtBfdQP
4ge8T426GE9h4DkOnHOQNoctIFhQ46dJi+dtCXw/luGzmuKa3miZMwDYyb1uzU3M
xaH8gZHZlIgjEEVg47FSB8/gWKlbfQzpc/4MvUnaO8YG8zNd32BQXX4e8byNP67I
GgCzllYe0nli5y7vWYb3iyMg0HhwDLW8MSbtLgU90E6S8MNp80/5FkbJdlHbtCrN
Wv+2aT7WyhMOfX1WQ2mH9Aedote0/UTr6scJ3dEySxDmIbwupq9ck++Yx3U7VYw6
hgpC9HwrcGrrZNy8h53ScIZjzu30vhB75yZew+bZEU8eHRLvp4ZbsziARiKdMLw9
psUNNyXy5Y1N3bN4FsCvAdoowAiPGZdZqNtM3oPokIDq9dQtisG4yiv8p6PDi8FU
6nWis+2IFVRe+OmeGSe6phzzU9HD/eRWG/fnXdbbqWKHGZjRc/TncODkE+o2rQ4J
cMDHKjDFJBwNsOOusZnU32L7kY8l2aclsMvvr7Iwc9Rzo6Gba7W+jdXE3kDqErdu
LjmKkkcENqf9Z0YIGXALh4RshCQFFBMCvkVl1eWhk1nkqngGBdxwQwhKtokB/NyL
WowEEMAZqB+Amq+jTSSXUcPkYY35lYo+vIEE3RZFBKsje0YiFLgqKA6tR4kfZypo
bGYu2osz4m8vcHnhZV3EI4opW0h7S68BnkxNX27/5XQX1dKd/MJ1ixVemMeMB/Q3
ywILeqTDnaFhv8FUGWlBc7/rK56VkpLnGtxRbXccfn24Zg9hy/jyKIgSu/uXzEle
XvLA/RybxHkfd5YStkCrq1JUWDoUYtKbSSE0/pj+VOd9CJznzpZW7b5NmZLPSxSa
e+elbugx6bG5/7yrEngUCMc190fLPnKclQybe0u5P0a2xbGBUjw4j9RPb8ZfrgMo
1rwusXXUKgsMa/MGjH7U+sRTY2xUePDCnuyX7VtpRBcDjm+DRXQW/kDNju+F7tqO
zZM8Nq2m7UVos6tko48R6brbDcEXG1EYlxK57jKIgyXFUS8x98EyLEXYcci2m0dh
7sl6SfdyPiuqdh0NnQkPbvDHIKvaanyohCpYAvvYQxsH2LotQfcUUF66dDAqYy/r
rOWpDsZsm8N6vRHwp5ht2bQ5Xbr+z/J0bC+TPmsazB59P12QNGI6wbXYSJCQGb1B
avknUA4g2V3mFIB4eXFEcvZdBq8tKSMZKHJLBgX8Cvfh618PnnISRXXPELapJstP
JcgEDH6xf/ZxI0WPt+j+4J2A+PJvGczTIgJeToh2yUh4xmcrcT+bURT53Iy2aECX
1zzSqhUGG2bs2Y2mW50uN/kLyCuqsqcxiIt15EtYcc+fIFNr9pC2dArN4187GQ5P
GbuNX0weqHpki8c/7Dxo0D2qtwEDtLsITifz7k/Y3vQ+eOYxaOaajGnN+G7Ei1aF
MGYdLxpFDAIwPtrvTMXxNEsP3OmNeQLZB9RguX/E7Ycr+Ombh9fOqDPh54ufWIu4
Bdq6DwtTSrPYYnXvi+JGGYInepN2aW5q8KtvjD0Hjbqj8MDuHXGPlbvpogffFOZ6
KPm5joVhf89bCbCwLL9n5BzWstCNa/ocuccmpKN8woFz2SqKskD1a5TMmdcjA1Yw
z4+OpxyYU2vdpk4jLlH2s76QVloIg/tcVTrkgjykUY8IYFkRYXHKyyeaA96Dnw7O
xSO/WhmT5lYCLjcbBlkCmfsivr96TxDmXXQ8v9ke+9RACeKo2YszjhOYS5Z0rg/a
Tcsud8xCftVxxV/ov3GKihqL+EGaskcFMA8XvOrKD05/B+DseKJK5nttftGWD8gZ
FhufwliQZCBYwZXEtzILLBonnRnQSbCs1/BclNjchvYddzSlOeBRigaGfaJ6EbSX
toVvhv0ozNwZQgTR8xYEw26W4j5zKPjIhifvXO8i63zgSEGuRijAN2nGZYBf5d+2
AzeDOA3kKflDrY2JhOw2LqMjaMCbnYF4D99b6WlE0fd3HbbeSXcc1P73t3x0y6xd
kfhCaHw6EyzhxFi1MEnk+VA3uDbfPwFkh0xUhUpFF7xqeGSXXZPp4GovzjjmgiaK
tcsJX+yynpdYhEUtJQL3PjwU5OyfL7TwDysLjQcdzPriy82H4PihqgvknSPehSdE
+OygFZMXUBmYouCxjHJ/X+SKfTkvxkDOh/mlfm3cWPtsKfq+pYK01Wd8HI8BLIKV
VrAxIq1BeBn/HGu1Yh8tmQDsGdHGEAJ2IUJBEvHQOHzyR4vq6wonlKw12bGTt+xL
xlA7sHOx476/fWVUWo0ELrDsSwqTdKmUMyeVK9L8/Y5WDltyaa4fruOhdyAlw8Wp
G0n0WcbyXtgENPr3OgDrrzbTNcPuAdIBaLPn/C6PpgKbrCOat/jPYU9OHqBfDE/e
WdlPr1GQGLYT8uOEaJWDqd33GaWr+6PZCvan2paL4VXCANuZ8nPRZfGU/Kqt/HIx
zu6fWCgh50L2jAWB5ydPNBj7fmUModyW4moqoYgrrRbZ6dIeKBKB3mQ8lqLcEd99
v04SR5uZU8aDgapUVJrVSwrpAhrJ33XM6yRQsnTCc8KooPcPmpEwuotbhMrH2kM8
nxYhUfwCwnS9gr+8INPttyjhNmIjvG7eYHJ7wPO1R2yfQ5d1JN+PNaTfDJ5cgeIu
eJdsnB8bjPw/hLta6gbf9/aO/EEShNL7MhJlAp84tDBh9KdfyxZdne+eIRYVFvtV
IqyW4eTVE/05Lilq9DF0VFEjJ2ixJNefAH4uD2PLy8w3DSKrvN3i05kibort7BJD
8mDn5qhuqUcLhshLYm3aheTbef2bqqaPf23RjYtxBoKe16+BJ3PIRkbairobZp78
U6pZWhbPPlliaH8hSTKz5VCQa05KZ9eVPLTluOdlWvUJZ5SGTYLwoQ6XUZbu3Eds
fE5xHV37xmSODwGeNTVQUtlhtONwdAQ1bSQmV8yeI3X7HQCF7y23VqrRHQ5btn7T
kd54pGLBa/BRtlUeTO7qt2kU2eN9jnDH3QJfkR15xyRHxBa2lLKFleJSH+vxuPv3
et2m/Y6cCqQbnloXHz5KTIqetgJwiDz8jS4p0k/5OIXWXXakH3edTWkkhJNezcZJ
KebZgjqccsqd/R8jjQnLiyC+YFyNRUdrnvZZnG9gNweeoCzcTnbB64ouf7eRbT7G
AqWC+/skTEVjhrjKrfbgAuXdbVS3RqetwwWhfDHYVKvZKmJc7Y1DPj4jUoVUTHdM
kb8H2OvCB9fIKaylDi+O1NaDi3ggr0r+1DJJUDQiRNMw2vgs+UK4+ynrvkYoCiTL
2raZ0C1HKwYBemJ6VNPewOuoMVuCCYQVD0GFHFWxfaeo363dT6HvUOfM6kWUvNVw
pnxzHywjJodZvT8/Uwh5/khLudvMAc9YQ0UfpFriW4GcCn6yf4v4LCxECMvuZSn7
CJEuoxnMRMYHMVDug+YLJlpzO8LrzHp9z43hsGCGNALZR+B6mJ1cRAvlGRjEi5+u
ZP9Xm39d6thYcvIm4nlxEMvyVES2aRuhmlyt05Kz8c5l6pbtIFPINNB6gxAWJmuC
63caMR/W7V11c57i7tQe/RqhJFJqyLCtBYY1SkPPz48e3UbT1crET8uhq+PqRAjj
dORY3H4MeaPEYiICm4GvECDX71PV/ESW5B+P4In+ystqenBfDp9TvAnZwfETuZh7
TJHm66MyYCGeikupE7Is95lpdFhSiODxYjY6OuMD2B/XEDMypKEdxYSzWtr4V9Qg
gOTGqRYMLY34OloRF4PXZAlDVU1duGnogTQC7ZZhmbGnUzZ919VBoJlgfieVrcl7
k4n/StrsL71LGHH/TrPZpg4Rc3lZad0m2jG3+DcBhuy8HilKfvq6yDZjWs1kdWpw
BK9Woh4KqWm72ziZmwtClmg6LvAdPVCiLEyxb/BkKM70j0PLb/DwkqsL5HGD8Aro
P98RI3eBekCxspV5KayBAB0TPu4oMb7raymuRacZYy/ZHvw8Yc1mA4RdvkgWdHlc
RvYoQHxOVpYXa7v4j/W8QhHCpxi0fK7KuEENEfrcCLKFQ6eBPbYglubEKccw6ZD1
Ld/10+frBD3fYc9uMHD/IaxiA3+gAlVwpFnWxuph51OaBg95x28dpZSVDKYmKonA
Wdf4kV9QcyhaAuflh7uJ7yFvUMxhRuKvazphj54O2E0c7OYvXQAalocuvDa6o+uo
a9mvvexaIx6neP77GSpB5tsIqQtNUTs+Z8iTEcY5A56Sa1vpB60vfU9165lwO9bw
ftVSWlpoxtn5Ikynrpv7k3XdO9UqoYkpZ99OlAg8sB5iPEMz0frjlv8meMXMmAWe
BUjtbOE7pfa6kPhXkViRrf5djf1jEiAJkW3S1gQVwmKWMi8ylJwUIJXLLrxXK5rb
eLdikjg64h1QzOmA9UKwMRyJ9mfDteawORP6YGlQvXoXUZQblMlY9mfq0tsnKHky
gnCfrXmgAa6EipQ+VROuCnRhls84e/zOWfettuL6lpS4zmBacGWR3HivBp5qv2ay
IsI6bcCSIYpavRZV5sS399c58x+qnLg1O4Z5iThZln3ckKnmWDZzjBTBk1hn4nyf
xsC7zKkJpKmBAbghAk/01vT5xIsMQyjw59GmYYxTCb2+KncrIt8FVV/Mznnsh8h5
k6r0NKV10OYkeN4ATu35Vj7rwpgILKYDMtAPQV8JZM2lg1mYnA6bOz1yQZ96YHcx
I9zu+cRY9RkVg8Wxd6VGYfiQpT+p72f291RaAddl2+7A+SBjiC347EeGjd1SbAIC
hS27+7oYeX8XHgGMoVDIUJrFvNNR56JOYK24+eCB1j0wkAZqMpohJjhYPUeX0k8L
NgiPlNrfFPPG+zNWa/YLIh6Q8/W0ylA3uLHcs9SDv9DVntspyApsb9t4j2pfKWST
Ey8717pK7pSDnZgDcDGE+rME+b+apDROfkVzTYA49UZ4MKo4PCXGirYjFtwjRbc0
QqSLKw8FCCjAp/226ej+Pnd1lyekRJyIB09KXVPwMYDuZNQ/3Df800gtnVOE8jwh
r36pArZSB+7LjBgOfC9C8Eriey4Ut+KIuNRyGfY8ppfhzeIV0L8em+NLqiWKJiVY
4tQGIMx98MZ1cPYQJXv/N0pWvibV6MVwR060JmYk49hpB5AbAr0QAP+0Fvm1oYU5
bqxMizGrU2qhktRIUQo3WZ6+3ONKacKvgOabc+LmLP73QjsnjFBVXaOZx0kBz9lc
fUUVQyyC4evo+NuvSrFuueARaiZOjc2vcxszZGbjcjF+rf1bdky0G+2xn0dl64Kh
80w+L6dPWGndbZZERZYAesxJjzcjXZFryN0Q3q5Hkzs+QePVIAw/vlJvXpxUkgp3
y0p9ii2OsxDOReOEgRz0VN3KDLCHov5lF2DoaPuBCzD4uu1LlJf8gh7ftK2KxDP8
wGsAAnOKpW+Wric22gPqHs8qW8WTcj1j8cg979X1QrQ1gOWMy/4Xwr/obHEzx+x2
Ap0K8roampYVqw3OuDRDNHn1aaU/ZC59c+p1QGSf4FuekwaK26HxcnRWV4Af3n+P
JuaKKDC1d++HEB+UqhAgFCWjfIP4Hc1REV57o9RdRiYV/X88HDXceVNNxXhjfbFe
tAYYL02o1ZeEZwj+3KfSXfkPexMrwFYFsANb/oUvqgEX8NxmcOIGn6hHgnDEv/68
A9cYITNSUR/Kkk9x6hnvMJDpchnCHXaFk9lHlw2XRImeDx/XzpyonTItBY9xizf1
NM/tkpwOiyyz7kpq+3OFFRExk2bLAYZ5/AUgOyvdh8BpXetrWALiRsUer6B6iM58
riiZHgKGmVopa+/tnAeN08aJOKicmlXvlaTc/b3vav54SRm/lFR8exNRxAxeD7xR
+2OglqcNxc8YJAvkcMO56CuMekESz6/SwN8zpZmk2R1H1/k1r1oZc4p1MSoePMY2
ngIKUVeyqmRB4oVkugQfgJnXp8G3/rGBgYUYR9TOFBCAJJXdEFuTRi2emgtSkGYS
hTFjyXNMH4bFkQGSYZuKDP38ZawLnnfDyJQsjZTcDH2bgEbh2dJfF+ENQq1GPweY
d1jpH9cqlY3dkWfr8ddm8Vh8pOWWMweZ2MVtu20XIn5d5Xtt7Svp+Gw1DiJKUOaF
+R1R4hqTyrwMdqjifFLLc79W4DcRWAI50I3Y33Elv6xRLhxIjX9i9fMnMY9IGBq/
Q2YGbG2Q6cidU7Uezo7k0bqm+9fdcDfWAiNyBgNcy5MiYJyFX7ZT3Mv02uMbfrlS
ZoFMJd2yijTxBsPbQPJtAb6af1BrVTSfnq33+Zz8DnJpjoOl8h51fuNfx1uEE2zc
hcrLglxdSviBkL1W4zCId0eQFXFC455KgvU2vVFo5c9WN+exKpjQfjggyBUvyg2x
qa9GclupLw2q3fZ2rqU1fWuuhmtq/MJyGhyZJ3vEUwIOmqwxuzyesVELyd8NKBX4
rhBzaa+pTR2Udbbw/nnI14YybVW2wF2xdFOQa7cSOO09sJTEAKHOPwCSdgvZN877
vfRgmPGrN52fV07+rqo7Lv34nsrXqLEB+D9cNWgllgB1vE01+GAW2tQLIwi/PaHc
IpdEm8eMmMQCOUeiQfGvVBH5REKDrIjDo0Im6h0yc/77t8lGul77hmXEslTB44qH
9aIMn2y4QL2htTl6jTeYUmOTJLN1Pzu6sBzJ68w5WmHnvM7SA4fk0BksvfurYdPj
AFYiCwap2J0dTQmfhCs3u4QE/rFjZdDG3Feu7rzjN1O4yhCJLe94RKkgYUJQyPUr
E7Xs1bZHOz6BC6t80qWJhI4wgHGiDO2iH7Tv658Z+Luadydys5wm1MNEPqlrEHe5
WBVyMuYpMPmuGl8Fl2TyMl+3p7aStoyx9FYfTb2mEiZyxC3j+XOWgtPhYXqB5tIO
BY5+D3Z0Gx6Sw+qAILbJo+SJa+Jomrjk/qYs91+annNZX8XO9zNReWmUlVkQZADk
AYoNGLIqQt+XlMwY41WJzIYCBak9QEDjenBFzjgkxuEllTm8fbZNo1ubJ4Hkllg6
5kOOy3YkbnkmYwljFA0Y1WxyeeM9Pj15uscOnfx6EVJlbiKXA+bXyxy3cbLN81l+
/LHhKpVF7nkggz4t6GaC3yBM+ziqUYOQI4Rdz0H6lTxxBnC0nEZ6f0kWjVzBeYNu
VUU9lCn2O+VddDGZZ0ObXUTbdXZliVrKZ2VtIo3XZ7iHQJBUuoj8OWvFlHPqOSA0
gHIw0riXIJUyw5EVnGrDHyYF9i96JysKkplh8+vwv8L+o2U+JLFLH136UswhX3Nx
ocg2luhW4qE9SHbU5tQfE/7EzSgDZTMJMj/d3Yh7RJOeiITDwGN2tORLIMSltw26
t/QBmpWhvQAybtmwAK7za4JPA76Xm5UjNslNBmnPJlk7PHz+2fVCaKwsv/AGBpfj
qXmb5ZB4zHFv5NFRqNNSKSvtg0RNsPl2tUjehV17LncEb2Ck6CbuPn0D/lqnE63v
9fgXb3vsYdNucFiY672mR2eye8+K6p2WpPTeyxIRyTMDYHgtGOavWRAdpzT1lu7F
mw9R6m7lBYXee8zIzO/QLq8B21GLHUFu7GWPE11Pji1yjqHZLVoM3d6bwqxzbKi1
YKKkEUcXg0sjarglaA1pJ8ca+YJF4+667jFNxcEYi1XacEAxFkFSWopoMcyNt/sV
SmRI5QF/+z/1OUHtBOU17rf3EjqF0yXj3veZccO2T29iIDP8hn8mDhRTklbEQ6T7
oLicjjertBWMRkYJQMZvhVqGNHaB7pzzA7JBLAaSCdPS9VjESwzxZ1CmBo0R9uxV
IvNAAyGwJ1ncohbslPFPk3tg0lk3MDgZLZQH5YZEhikeXwnKjbN4bt/IZNodivwG
14MrF3/S/lbaSQXx8MGRailORSMQ1LUbytUkLnayBOPRtP+6INqLynbGcaHDbKGj
PnA0tQzBlB1yJuXGywYLi3zutTh7euuA5CVnHiejwnsFVuXceZKk1FiFxPyF3mZX
9E/bL5ehW8hZxdTkSFaouIz7fE0gGVJ+WGnIizw66r9Ph9l8gOGB6a0nvl97D3qu
3BI01ZspjD/H4a/PNUJDfZQ6Xsh0nj5Kpud/eKRt6EQ81+3dPO8EESZcOvIGZLtH
ApbAz9NWk9XcAE9nF77pf+d9rR5tdBng0eRwYuoNjtIO9q/fp5anOG3M7KGsfEQO
j3ttFeZBx8IAoSiCZ/uTu0H5Z8Lb8QRWxQM6j9T4tQ49+jVifkGhc7clbMD2xkAW
b7nqalishp+LsFkGhMwsn/w6FzQ+KCmapOgD5NitpAoryx4F+UTzuEvJJbqaGbFq
mBhN3p9atGU3Y3h1NA5S55FbwHLAffOdVckzB2eKT/07H7zERP1WyV/dBQ4Yi2um
LX0D9oUfG4J6K46kVgaHJWpN4k5jqWailXJm/Ta3zWuq7v5LDuBVLODpy1z8Wv9a
5Im/FXUi2zNHBJvIeyCzbf3hShDvkhxIe2puA51ez1T+0I5wfHEy6CgtEGWQSaPE
XvBD0LyGVPOX17nxFNS2L+zy6Hj2CkKFtBbG1bNRHUaEsh/yeMd+PIspYLcD1M1O
6ZGrdRchULbcUY/xGxWgL5vfbBfmw4ytf2I2xHQutLmkmztPPkYJ4ooYHxocQAWq
BIkyucQAropcaugwwkWX4qxwPsJiDW3B/GQI5/sae10KsP7geoc0pHN5limrCl8+
T6236jJRFmQ0PKPwomPK7B4bxiUYlob4RotdgVI8cPgBFUFyagPqYC9I06tfzC3R
9XPlYPWmpyth9Sjv4O4lHbuz4xNpDBkJsK3RTrMSVDDwt0y8PxTeESPCYv7ngIwz
iyN6U4jk7Dt7Y3GOFXQ5bNQ2uOqvvqEPAItPp9NCLPX03On9H4daqJvpTBD1VcF2
VB2j0AbpNQdZX8ux3tCsHAuP6WBplhETrrPYUHzAfZ4qrBJCTeMPSz4BWR/TBKg3
MpfI/Ut/qreMugpDKB6CmO0+yJcK5MeJIiUw4Nq0RmDXZx+3joF71JrrbXxA4sAg
4FThOedSqEv98bHW8qy5BU8ojCf+6Cj2kBigIhTXA+k9cwreRxLlWvxEWvDioGdK
UGEN7iVqEOvBm0TzeKjf1BpG0LlMoAh0nmhFwNXx9il/EaUlFDL/pxMokIY18pKr
XTdFMLEITfjkaYNrLK8+YX8fl5KebUAhWrRm/E3fpOKoPX67mxvqFbT/xjtlfCYL
1L8imOXCU9RDZp1DbvXsf0WpyCC1oq9pl1Wr7lK846ejwsYHeQJRQBBCk36hJANp
VqSPe4Qr//SB9kl3br6xo69BD25T6I3gLnckNbkP2iZeuj6E3wt3i9CXPDXhTFWR
wgg7aANyK3tBe4K0NdPgVKhySV5RpybOFBqLOkAO9hZbSomhs+EZfEEyfVrmPbwG
gQ51mu81jiBSR77+zM6/rHxGLaD9+uclgHwb3hdmG+yz+AawKWeSIZuIJ4b21Vu/
IcN85j499p05twar8N7cS1Be/53HWB1wXjuwgLgcgJcEJVdZP1ggIefPcVAix6y4
a2CMHNYKWiJ3z5bbUpP9+oBVt1LCwJxUxXWg8KNIluFOaFbjGCOZ12cqEqzjPP1K
RRKXcObYtGPZDf6MaSA++nV/Sh1mCqo/D59CIyPinCfPRMVRfzKIuH0ZcqP2wzG3
tcW7ZBlVhFB0UoPyrD8WznZr4nXMmCK1JFDcg1slP/njidYJ+uEOJ87cr/FfsGr1
eCSfC7BEX7SJFz8W2unFUqofFAZdCj6aR5Opg0GGcAukkpZdoOnNE+3adyeAavmk
X5L95FN7cUjNtV832ouAu24Lw+iamqZaRpS8HkyAjneyzgo1rOhaw2J1wwHeF+PE
XWgon3b4FHpxihRM72kiDhwtdRcmwJLN8pAgPgfsL+hfmpLYh+qhEJ+lZ7K3V+3x
q4Fm57DdGpmG+vk0n4AywOUzVnxths3qrBYWrFQ6rpkJbhTVCwRUKpQMDb3Nanep
OUXoVFhxnf5Xw1pdNWUnrg+b623t3SFwl0tGPYMYXtVxMMDCgJtYiXAh4TZVydjw
GkclrYj4ojH5PKbBtH/aWlhMB1Bu4Qk9wg95GgSxRS9BY6muwvjMki/7OG6dPjup
Ht86X/jPNeqyqgdLbg5I9PNeiMmFT4QTp3MxJAwxBz6JuS7ygIAOpKMm+wnoQ/Iz
0ZISDiAh0wqfgMETPEtaAgqy22YwgJfNq2WgZuYfGVTxwZPwXVwp5h8CqMwkxosK
iC0/WQ3eRYYYfZnUwE4tmnXepiEtJUjHj+3QcQw02OeHVLqC/8ewAjfQhgd71IUJ
jzprMsyZBxowVKuMeKlGjJN3rTjnTCkfw3JQoFYk5PW6GnQVTYQs0w8CWNmJYvKG
zylimJV8eOm/Ofl82bCKkgJefed4oaS2XwuNE60iwIDkDE0Ac9u82dg/GMyKaxSg
Ptd7KmZSMQlC40ZUnbVV4j4AaCO831vUmkWdoXn5jyM3iMdtDOYiflMyWSkpq8nW
UlHSEQzkh6Wok7eoIPHH1vCMX3dsZEq9ircVL2pH7D1XXriWhlwxVATCW7lLsW9i
nMZdXkZvgcOZmPQGHipHcDCleZdPf+YWagpPB2TzZuVXhf2wczwbFAQ/vRfPgFEK
RwEgcnvp/pSQ2faG/PdGLiVsLMWkKSPQiw33r95KJ4KzKeZyYjX91PE4GFOd5usn
AzSLAtBymS43FRhCQFgza6VtAAbv2MdhEoM8bvlsK2aKxrHXu6KA0a95h8tlfj22
wGnZP945MT81+ctSH4svvhqjO8Lb/uapkuNV1lu1P1DqEJaU3OM96Hy+aku4rFK9
OLNggNAxyfNozboigera/W7SQ/2FeA/1tuZYXUCI9TIsJFhtAyuzSoMOe2KKIMoE
PSameAjD2nf90HtahVZ30y0hDWaHtDPaooAwlQW4yRhcL1zvaVjmk/38MBf+A6uY
1A4BSyTwLGL8HWuCty87Ay/mBA5RjZLG7Ca3X8OltAxSzFtePzom8RvyhqD2CRSh
RPUovurJdULjgOHOBUVRuPVOqMW8HRnshBMEVM6oNzl016r8HwLWVKqWqnPNxZjj
jwfmcSmdf7gmp/l9gQKnl4v5a4MEBYf2yBEoKFqBn/91/XgxxBzS31FWTg/xW6TS
ojTKNX9S5fSMjRpFbAZsNjmWclME+rUc+FIRsrPlK2Cas9CEhK2hwSX144cWE/N8
I6oEx9ZyKl76uWIbhpm6KunrCXRRpNGFhOZ/uWwn/8CrHU+qsHJemkK8rUIzhxBn
V7FbQ6RuinUvsJOrn+c1VIuvLtfXwZsjEZpdTDBlVR4Te1VvJ7nv6Lj3UEiLhiP6
X42pjVvT09wrKIA91DIO2S2395rcwt0CLeZBL1d6SEy7+4QCrBE1WV0tSWjy6sAv
cwtrh8bRAk19MDvFABNR0GyOYHg3aHG4D68h/Uk1anFjU3f9IzJrzaJQDEKy7lc8
tkT5ltjz5PpitPu8YG+8lwGMHEv5gImqpnLzWIinAyYR83fHw4MgM0Es5WJSXgEE
PlqfkRw+PZZe8CBDsfOIXrC6cNlj9HgghQaYrHFeDN1SS4dtQkx9dabuaCS3Zr30
kpETwqZ0CEQXRsx9Hbt7CtXz0PHZbGiB1K03ltvDNDqqoRm1PNhTCxdHg/+obe9b
JvMNz+pJg6SjBa85+I1OLDDSFW4fb6Li/9AuJWFPDKZf1bmkw8AtSWKZgtNOr1Qo
wxQlDfkjbcquSqnpUxMgf4ahONVd9Lz/wInkNtfIUYKqQGe14+8qID6k/m0PGbmx
ERcTXQosGAlTaMoMZPYvnlSolip9JUfAGYC3Ca9lQtHVB8eR32eK2HF65Q1krQxk
LiV4W6OPJyAaZft5WEN5OkW3ELhqQ4a6LwL2BfGzz55fbNuJbq/+i0nJYGslYBIz
BQym3BfEQo/SnYsUeephUYS8IUBb6/98Qd1WiiQhOuQbKL4dN2AUMyx6fRgH6kJu
L/e/QwPJ7AlPghE8Nvtwe/Py6+D15u272ZQR3+tuyqD9KZBZGlQYyivBixCaUu3+
Aah2tpMIzttiZuFhbDleaJ1jXKlbBSV4V1cHVT6X4CEZ+hGxt2QpvnHpm1TbUCv2
MHrsAYKZRl8OwDVe6/ig/KExUSobnxSvPXddETW3Oiy3dbcac6orVizFQnJDEejv
b0tHXF1mjHoQIuZdec/nSc9S1c49nA8pFbelhFRqO89I8W05XEXKC3D5bmdh5A+R
BqXAMPHORJt1CEqjSqKOjtK+e5bt8+EyhdCAbCSsXrAM4IDYfTLuvo/NzN6sbI24
lB4kM9cO6Nhcz3JbkcbqYKMRA4LMHbihSRZunh4iUKRyErpGFEMNYsOcdOIHiMI9
dQdsCEiH0/lDvL1AgEw8+C5ZCun+U5EM1FwLjI3Kr5AnVdKBCEK5fvz6EGwG+xDX
Ecqzhr3cBMVGt0BgM93LAukJ9JcoH0Ujlcm1NcghgivtY4u9v7/1HF3vJAbRdluT
zZv8ld+FYwr7BNF17JQMkgIGMlniuKa2VHgS15UEhZCqwYpfUzNvY9JpLLkb8dPM
RAjLUNpK5x+XWgnOv96VOUaw2tGklBLO2FgsK0Hza5v0Ja2BjtBZ8KJBUBvM/8QM
43k+ZZy51ZXueKF2YjFlVX3WAzzje6dR2otQw7irlP9lK2IK3QchEQYqQn4vidvp
m8wrfDTSQMWkjAFcTae1VRqHUFve8t+W9oIljPEkgU9NBjm+8PoumQY4mjWEO4Bg
qjIH9pzHgUpuFkAEZQ7fX2Vu7r6G2fnKWQT0OyWJvdTxyAUvzA8ttpjRDLbayOaE
34YAIGwBgN9WnDhRhAV2kfTxh5m61E7gqtPNZBmW2oNS1YvZREUPGiDtmjZRWz+t
pQ6gTTb0oKgVKnLGEabfO7Nyy8MowV/A1SMwK2PK9i2bd0Jy8mI7Q+ba6jUqZdh8
7Qk5gRP8nCi5llJr0pHEzg8n0snZkGrXeRsQVfIumeOIZvjuH3QX4WRTWyQ98/aH
7pjG+4clLKBqkfhNkz8Z0/tQc2wWEX5gX3JqzyDdLFSi8t+9jTgg/7Ha28YoUfhf
G7Nu3AoyLUUTt+Nkm/eg8Udw7kRSP8l7lGwRwUltGXhgPfdH21h/lKDJvR3UhC8j
auuc19wEGGL3i4WbyZZkrPD01ki+jmn1/+XELQhaEL067qvjfc3XQOGMVJCvDhvl
z+lyIX7b5qWvAZxzs3gr/as+CyfKFerxQuh/T0+QIF0qqfwdeo0vBiow4d6sDQiw
4NyHZ4iKkslhUKlmTpoq984WnqKUcyRQVI45ihYxBtANawVCS/us3utTxGah420y
HxkbA3NwVa0IdHofkEhNwm1xTUBczKdjFePgl7Kaf2QJEcn4DWMPv29xf3Yx2Lwj
jCi5QfM0u+NojwYvv6o8+SFzyT7pW0aj4bVQ+6hnzPc+csk2PqBM0jngb0nNtGyI
W6OJXqE1QLfOj7VrcT5LmU7I7JIE2hyF+vGXGd/QiQmS3s22YlGWn1v5gEx2fxT1
Y1ErQone1haSfzndq6O8Z6TfNTbPFwpfYqCV7JI+S2Ao7mozBtS5iyHBH7+x0mCO
qBWG9iW23fYA3v64/pcvfAV+3X7pzh7Fqcz7iLg5B7Jm6+5XJ0miGiAinCvb9VpY
crvoBSAEIgYjRRWgWzIYTIPkmMIqRezcPC7bpkzHeQbVipMJKpYlo3BSVpb7eGFw
4FHgQWHxuowTMn/QWV/ECoY3aneMu9AvBuEu6L2sxsns5LLuXxcIuSCrjm+jpvfG
ZdATkFohoi1vtGRBpydWzoiO/dBnF7dgg8jQuEorYo52itYhM7gIljG7OM0n/yMH
ytTFRtap180B3fluByDkm1yJNKR8gawohWP3j0rUtnomHELmgnfOPkU3HGVaxbcX
tushjE2FOurc/Zc672SElj6Ktu2gDjot9rNyCT5RVHpe1xN/txwDjwKOpwQ93hgN
V52iWvGz5bbb0bC6g91lI2c1sjhOXmrBF6cEaGMxUIqlxyX/mWhdORlyNTSKr22V
8NmVy6zv40aKw2OxZ1xl0nqULMEJCGukUZwzgQVS/NWMebD7zJj5A+D5jqLlnviy
svWNzjOfFb/Q7UrdRMsvL+GJyaAgHtDGChmNCcXTbP+rXH4q6YlT7KPnUXHAu62K
BtIKjxeniRq9Q5f37EOF4XKkx/RTTCNoEq+JRdyBYPY8S6ItitKkPhD2BuSv0gzG
RFlNyyX+KTCTimtOpY+EBLJnQd/wGkVJe6XbOUIDzrU1TXgqR6Ylgr0ZRkDB3DRF
4cMMAMi3vsnSqc75SqZKSxe6fx4aJsYEnD8uYE2kn6moOY5b8aUQm+G70gEI7Qfj
rvZp2yXbVR6o/vnrzU+rN5X7IkKujWn8qNX+EgDxNd1E9MB98RJ7wIn1qQVbwEPD
MozW4OUYOQmRAjjt/2TQj2IlSbcLJnwVk8Vk23Wu+pxkXWpNqxxIpQq9CT8Vm2KO
a2UmU6iQ2qGDpCvK6lAaLSTJN3EuxF1GSYpXV6WTDV+GrYXoI8pgqbYpRcsm7h+9
ozjerf1yLMIKS0IGWmt2IeuBFGv6Lz0jIfgftp1b2H1CfTDcBj+8+yzWbeN9KQ4Q
VQIBl872kbTxBdBfLi+DANp2yUGZaKEELkC0cPAKVWXSGp6sMlhQpkIC30prH52B
ADf2acvBUBKTt9DhajV68/7vr0CKut3+RaPmFs9wDMDVbltF+30hYCj76SPzSUEl
4To0B5kkmTnsvoBN9hmhD0h4+ut52wRpyb/z+X0dKdAtGQIoOzxsj1sOCwfJ8b/2
7w6Z5ChYU7/mcloUiOD987yWwFpxf//eWoeKcaImHG2nrIL/xsdBhpy6D4jZJCrj
7LjlaKEBvVH3cVIpWYadnL4PaWN9YvYsxf8dS0acHLyJ5ZZZbI2HfAoAl0xjo1GU
HMqRQ90HxWhhCjBmOHYRHwLKQuYLddAM0wpba09xA54Git+QO2MVWIyZIeWk32Xo
IHbBDtVvrH9mriS8pO5s6SLGXphQwkOnkr/a19ofgJ3eNBNvAwSGI9trWmjwatc2
j78Luts0ebeDlK+cRAcbFrXW62019T1jveSm+HWT5XUImgT3TqTbDhkglkJx3gbl
syZjkKmEPzPfVLlNv/GWB9soMOOXKqGgREMcVZCbXAvM710hRKL77na/TxBaUzet
k7kSO12I69bC8Qf0mTlS5oO2ZhGO2rQYUXM9ET8aFvEigqkHKzpL5M+BnW0ZN9H4
rWy1U0r4qNIEv9GLQeyfUcSUn+FwLCsG558anBeLR8xv+/rLrJbhr7jcfIccFok0
gEzLL2+ok9UnX0oAOw2RyCekuemElGw/vPcaPZafP248MGktNWlk8Bio1n/VXBbE
MEEQdIIn9mGz4cDlA9VE9tTlwICZahzOY24ugyeU4y/579yiu6BgdnoQFwWanZIs
SNxivP7Av1xVweuKKrnFKM+RcKwaWpKFhmRAUQBSlsY0mriFGxFRZCtB/0LcVxbE
C3DhvEgnqvMhwW1ubW2HTRAjjDrmnPOp7wHHgHc/ss13/KpdzZMUv9k8UoTLiWDO
5oPCPhao+GSR9lDkRAPMVRup0zsBX44T7dkWGimGzyVbFHYj7KOL9N2lxfbKWBdA
9aVhXe6RIT0VkDly79spy+OeMK6A57ju5vA9V+Q80YkLMiRDYdz9xSweqa5HdfD6
QCYKTpWPOS77gLhSoP2KPKoOqp7oJFJvVqvN33m0PVCSwsfT6O6teUtHvWRIH5So
WI/MCS1WKl77b8DFdSa8McfBSdnZAwq7JNJXLcI77tB0MShgRBxAJZs9Eh0X9fNL
lRqqC7UcRw1x2y908cgw8LZSrAuriMEAjfY8luORqBWuf3P7t1pQlomShMmt6pmP
6/flCfsMgXFu2UNG5lOUkKE+TR/boOh8lSNOndI6knntRdl3EwxIpvg73BOAclEL
otPzx+V9rQaUCJnhEn3jo5V4Le76POOWZkTt/bM9fnHTWAivWk0pM9nNevb+IpUX
/R/13+osb3CpfFoslT5E/8hWPxQIvPraIdgh7mPrV5gTTm5+7+gOPyk7nqOKjB7g
dwpBhg62I+DbrekmSUjJI0KlTh+8kavy3lmVU8/s2NIAIHoN/Q2YehIK8L5oElhr
yHsGznDwlPNTtfEFutb753HfPOnYjR394UQjg/frllYcU/vOsLMD1DnaFztK1gtt
5yiGLmbY+JF5abSHOHDN9mCYOuDG2XtnH/U2YLqLjqFjmcPBOSbeq1VCY1PyFSep
EXu0UvRiOS4w5d90HFjZTrvLoO5g/G34bH5TU34nzs+Xhmi2cApGIFbLKRbkKIxI
gxz2HIFvAyyb+yCYLDseARTJ8ZceRsQMfusmxXFprjA=
`pragma protect end_protected
