// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K1RrJPzFKHBXjasaInYsuD7j8KDnIQFJze2+vz5SlV3VeS3hMSkY9uZV0f6QlRxy
8kwegwSvCtdUtNfR0FUjcmCrCZmtYbpMVX/nQ9UVfQK5ltxMrCR9T8O/XP6fAJ+F
dFJi4J1RuufrQpVm4trmmDjpZl0m6b/4cYM+JLom9kc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9776)
teWqTQaClG+SCoIN5HZD0PJe/VvWT0BDEh+14rZoej7w2iK/s2X20uQtVJa7yxrl
jpnA8tO6wpv7FwIDVfEjlTsJwPNjmS0aVT1Vq0ARoQa3AHQdon4sv9NZMey316ku
q6AszO6aIXqaKa0ifuFO6luUSEXI1G7w0rRj1ZDdyNMTPHEZlMWnz3eMhkaJc+CS
8qNp4Bz+tcS0yYbhiIVFql38A7hqhsrYqaTqBuTyGlVSiwnhN1N3tXK4HBPYvxwy
LVh2Qmf82cWF40XS5YXfNKeeqbNYqPJ4+whGmenbeGln4XYtKTrbEtcgVheh4pXv
HHiyV1BsDPfnw4Ej4O55M15LGTgmIleFEUM87DZwH+ksUe780LUdiV4bvO7ZQDML
RDwWP7pgusoDvRsHJm+Yq6E5FJDlj/Hfg0xIE6DSBSXwfTdkEcYn1gFIDcFqkj5P
lnHrVz+PB5UaRYwfeH1Fh7vvOrYSyq3kMuJg3FpP4UI9E+liRIWY4hugMRsOpqhr
5ZE3tx/C5H38ZmaGZnv8JQZAvS65QYwLjhUARj+fk4m/xSxf/A70YjFLWkoXlVXO
w1UHT20vpSknzY/bxhlY1loaiRJ1SuoJg0+nQErmgZ/1AELF8UzIj48PjAqlagBF
D2BK5/Yc3SkZRy2TEnzJ/Z5OW3upndOXWdj0g3KZT9uNr4HtBa71JFQtifFC//SG
2bLS2CH1mToPHC0Vhthj83zuGeu6FgGh+LovjuwIYi//zt7PMeRCzEbRTPA3PmPt
rJkLThlSkHk7kFk8+oRTm5ravmCF/WtXR7gv8yvNH4lXebkv7FrXXEsR5Dqzlr6y
cgYfuHkpmg8rwtodhA8RFdNrc0dAD+FRCqLUMIcVk/5IU6/UGII2NTNCD2rOYiR4
/c41jLCXyDW6HF/IP6MoiobM3ODVcnMH7ZCDhK9GiCKSmThG0XbM6kb9Xv8H1vc/
7HR1qkGHjFtmT+mb0XRJAoWUci4wWM2Uh2FWEr71k9DchurMWe6SJ3i9KI8bStt8
qIjP+Au5Cs427qDe8yG44bzD0wpSx6vMgMjNfnt3P+sJ6opFwMthdZb1euHjCvFK
fjxdVfS/ad0xb7+cmGFcg3c3EnscBUijw8RfOWXR161+z+yyAGCxTf4kuV05hjya
l4dCET3PKd23r+cCkp0lUQl+xVG3cjOODK8BtZfBHTE3tfClcycnMaY+TAna2ko1
cuI9SnvoqzMwu4l04dWO8cf2pS1E+0EhwlTDlakJZfak29VVHXrvpGJ0iJ2Iw70h
1KHcKSqd+MWpcUTSVjjNHmB4Ge4rgBOW1orUkEPlZwQE3t9niNz0mVFz5S/ciTHK
rwEo2NL//pzeNPrvWlh43drLYup10GyZUUnYQhr7oYgNy1aKELBoAkzyjR4DkWy/
BQQJxL9SyWyMb1mYQ2CPc8eWbgdxud2rEQ21O/t9Dr+I867Hq+1Fwg+AQtVbpU6T
nHCc7p6z7ZzNsWQ1o1upY3ttvZFJ8Zlb41PShEVTUkiTry4MY2KFmMB8P0JRT+LM
nJbaCzNkZ5P9FTNTHltKrrJFiQHiyoji7nn4EA/dby/TV7SZ0zaR0rnpOdXlmMHE
7SvrVcVDXh7embdOtb4DZDiE+9XtqfFhErLVmGlrp/igRBA0rju4+Xx/rkWeZDq1
0qlWvCr6brLxwEaFXlDpS/QAu2atf7AeHBkapcwmAWl6SrV7UhpIGZify2iBfXOD
XTILscOA5ydNEPhbOb6z4qa5EFDcHpXgAuQthZUEdw+WsV50V4RleH5oqvyR/9KT
3cAwFi7JLw7+af8Mn74s8uJEajWjrzAkXhfiGuEMVpisXnD/orarFQbmsw1G9cpw
NSVzBAP/6y6tIkJj6ttLqbOEuDTqcvy9gvNCkCph/nJwTpkuEkIFgyINg0gV8Vmv
ZQ3xhM7HUfVSGOwwnXHtqxFPcoUSip3izeXGlAv41eSyBE3xqRtS1n8gSFn5AUrq
hNshlVsLUXfykDwn3n4G5U1wruasIFIFPPCsnSj2jOlRqZj7WotToE4cQw/yG0x6
Z61955VSLiKK0ejTBmV7AQU5P8avsu+jg5x31dwn1W4iOYWloDrgf/z7es9y9+Zp
CzWszY5DsqTl/+Q6T579NeRVyOc/hBdom/Zq418uuKiz7qz0zwYVt0kqYPD9NxYk
+/w5szPwE1M7cdMD1HeD2P3H22PyiLQS+2zR0xk1DznCbjNvo3MsvG53iGXDYj7+
cxBhJmQs735mO8QMgmO+9bxsCrB0lMBSABkojvBQ9evBVb9JtInIxm6YnBsgN3K5
BsKk+yf+jwvtU6a8NPtWNnNESCbF0Zn1EjUY9UywZxFxF508dWaOpuB7fSB/8Rfv
1WnWsr+zomsqtY2DAyMuul7l2if6mDWLSY1ZPa66X/U0OcggtgOWebx1D7+D/VPw
2ffsrqupV5cQfp16WtTw3Dv8xn5AggdPOo2l28L83qeC7cIhwSKza0mf1EalrAXY
SrTkiqeRrAwxuSzQGNiY04do0mZ/1VpZfxEZ9aM/yduiM984F4oVgKTyO8UIimfX
QKjHorIE6Wjxohy82zcCZCqnJjOZNn6Dw7WE8yUgFdAIuto+j2YR6lVQrdMBeHSd
UAGozZ7RBgvyl+tuGy+Hk6xuZECrhHF0gnppVfO2FEEizo58FvzoGGY+5okQ7rvt
b4K9pBs4GDq2rdZbG1EBHZ+ZFDyFRTPCrMYaVkEjvrmJtHXpQNAJhvJLNaphLyJf
TNp5K5mMxwPbth0pamRSr9cRQGt9zIVlD0b2/1+7WRwbS47UHQ532MI/6+MqT7U5
nx2J4Hk+LJQrGsKuioeaiUc4l41BNm7Sb8v9FdUMsLeULcbVu5tqvBN5RvHPv4+2
uvaE/upNpObRPgHs67hpDrBDRAZzJrzQc/1SduxaWV9gtpy8WYetiHT14JxQZh7D
ZikWc5DqulGdL3hwHSYvLM01bojLggXgUX0depmbswAn548UNpnXJ5ECWlO/mPMH
PuQ3OIOJfc6wezdVyrIq1L3ATv0ysMYR8QIXp6QlTjNsUzwfpSnCtPmJEIYb46zR
IE4wzQ+MvIHltj9lqk/YhsMqCK2MoLOoKjOdnNmmnAkE+tjuzJIe03/JkHD/M1GW
ZPOaAfaxK/qNDy+Bpl214634ihnW6SYwXbzeh5t+IXa4SogJPc89iQXC+xjK7j39
ugvk3nVeJEEJ//qaG/un5Jm7LTXnXCeDBlej+5KiMkGH7z0rzcsOuGZuz0ZSV0Ie
g79NISHPjjj02Y6CXKqOgeOn+Th9BMqmol15ok/GbV4BVq/PWv70Jl2AOiF4k5BR
sb0zn1gRoZGyBc34feqQjaTF2l3QoB04YhUkvFiv3Hq25YkywuaksOj8ghm6Z5Dd
u9RfEF+VnAGoCxOQ1nKTxbSe+af5xexmaIlzEROzArRBDy0IsPs0sp1hPjVaB+Ay
w8lqNkOr8FWbJslop1dThAP7ch4YJurWyQMb1M2H6YI5mVtcJklQ0hVATHolVhLb
rKN4IZyfcRhPuHoboDP2mNpiFVYJz+cUHW/Zp8jmDtyu3M9vf2U8Erz0K6YQOaIZ
tcsm7IF1obVA8OiOKcUMQwRzkig1DwwUIWCyONPyoZqJfRWPLj6kqmNidRge5bJQ
XOW2TPHT3LXSa8fVcufiOBAiGOVctMzCPImveXtEsq+32yduooZTamkw7i/wwdFn
LFeeNnsVeH1fu+oWEyx9/hqJ8qAlLoNdFl4RMDqQimdZAMogr4fxBtk3sxIRoH4p
d/tofAOIxxeSZ1OkS+yvCowC52Vx3ooYWCb+6t/yk280jAE6VnaHF6PwdT/IZACa
gzIRkKEwQAaeKpqfhPxNcUNqfrHXP5W7OzmZdQZ+KhgIetjq2Ppb8HOKo6FBCWtY
t9je6J6dME5MwHMNNApY+l7i5Npw+SpCBNguwUfar9OPE1dGPgfyDiuUEGa68JeC
4m8ILZJVpTbCtXBRGRahMNQe+rAbdXmaLfFiH9VZH3RAYkZetAmBoU2e5pRH06r1
GsyuPzQsBM9QwTjiwoXoNCJ4EsvbtdDnjVBG4EyC0ybJXXd6LsYFazmsJsyoms5/
AIrmhn/b+gKp9RsdjtzJ3WCZKwZgyMihevTaVmFGglAVV4ZB3E5qRQ5/q0sOxQKT
1aHQDqybwnNjMg77cxu2Oa6I4CntPO1wFxVT5wogv7ylfs8GMAHm+V5mt0I2D+Li
o2gkSpSskdoMGL5KHo08Vxrxn09kxxIS1dNEXWK/91iTxxsCqdKNsvtzWzFdGf5x
UzBo6Vdrg4jrmzUvXpn6CtU2v4QsvZHmMLtdW2FwPLCFhg75WPPGe6JiB5UW1xs/
6O+BYrHkmwajz3Dq10VZasRF/wnza5VpduL8dbKiRXvS6/thk2V+2dPKV/ry5Lk1
mAjp7t5WtpHajzdfxbQdaP+42iHpCT6XULCzoR/NvkcmFK4oHHcRee7JP7v0SQOU
OcxQDPjJ17Z7/u6g7ko5vmNbPfmsWrVcBQA+araxeSVxTcOg2Zwa0ulRkyhUynW9
/VHeCj10CLfGMQ/KGaE56vqLCA/ernWTvT+MoHfDrQNRfhabi1WRgjb/jdoUngXT
soIA6T1TctFSMY2uCJtcnFSvLACUaC8vupJPP9op9+BnLMRie2Mece52lV3YF+mt
DMguBsTBe0kofO3lHTicfUHArasrc846PYuK59OKcsM6D6IF3p064YjHtHHb8sUX
MdvJCC+65aBqYs67jZED8e1sJCKnWpRx6mIFrChzjNzWwSDh70occQLIWAj32WTO
MObYZzYdQ0N03Sz+LPOCU+h7a5fhYpZ/FtmByXlnIkQgERAJkt8DmaSC84dWNhx0
WWtO8LD9WDKPeVUU/naxJtdvJMclHvn8B4i6JYzpSjPJktGvaNXiuUp1nhLfw4KQ
8Zu6+wbhiNvdtbBkplF/sbLKhCslfzeRExcUa50qMivxiGQ2KBmJTD4CPFuCQT2p
pJO/r5iw++nuULOzz3eSpBnJBnEoBg5mNeaUIgUScxWCgXG61hbLrkwruM2Z9wfY
QFcK0wtRJUeouG5rVTsXTiS8/wHsQGOR0XRK6/X0W3CVefVLgEYXvhV7GzEGPHQl
xSNXIqvjoYzGmyO1/Lahfkzc43DINL7PP3mK9KbcNoiyvGFRPYR6kz/uBFt0Iuwd
Mx8QqQ1dHFEgs75NtizQF/YJ2pqih+7yPy4b9or/fxDLBchqB/UvhiqLRne82c8C
KNq9jskVdIqRXnYIYOiZiiTAtC3NEuYj8JrHl8fYQB3cHVVUAT3XReAojgNaxky0
kCjWagCPs9cCtZS71+zf8qKsNXpA2rEZ6YKZvte4vDOdyda//SSwKqjVh7wIPEVf
j5uYjHdc9Sus5oS2oML5sE30mqi0197T/JBQKZUXWWvFTRmhk+P7p4aaDSEwb8p/
+KRCWI6wsU5AfrRGITvCRh4fVQ9/SRRhZ7mLSnD/SSTmoulP76YnL/0YHolaXND/
Ah5X9VtyKrlUEjwRS/QTexC5lLL2TwCl+tyMwaxUTUV+aZcmIsW0ungqWy8rTGl8
+i0VHahkqHm18OxLT2jQl3R3esNRV1KA/3E8TxfKyoTv0EyF7C1pjBHr0GV4YoT/
m9eq6htIW1XRxLvx5Se18gOZXRWD3hlhAD7tizcKGImTWc1M3r3vQfPEjyJAiCQ+
pU6NSjMlPjp2/bSxNEgnhtiSCIG6w6XM8CytDUnklihsFshAIGsCos3JOMHeF0TC
NYkVDbKJzfYOMUSPrVW+j/MH8mivuU5AMKPTkkJQWSRBsi90ecZ3/OkLD2xBIftf
1i0gZZpSRrFRXq6gF+ZIa1llCRNCQ9v00SdfGOdX1jgt1odLD1X1AHfil0Live4c
XtiUwqjLcB1LlxyJqO4/+6iteWu5+j+etbd+aJ2Qx3fy+a8ceYpE7HWYHyPd+liJ
g41oDj3KIoGPQzjNZiyNZsGXXnD/zepsvb70IE/NWWZAhR9Wt5Te9YXbEZvI9PQn
zG3X8tgKpuZVgSnwi99ML8zYVAeLtpzKhHTXJn9FKqY+GsFSSnqcSqnCKplNfFAH
RCM62GvpLnG0+qdjLYHDrH1C32jfLiBbnPvC7dJyiblMNX5CCmbkIF5NJlMj+MwX
Wsn57HsGe5oF71ozMorbtfZz0F61FEqmBbxiwTp08wLb0HwmrzRVM1tIBtyJeuhh
ILlsCqQMycjXgzrBgL239O9oqqfCtD4k3X4r8YkHPD0TFbYvTcV9dmdGhGJw2H/c
oMEtthxROWxt4UztIbnEQ6HSCr+N//g80E4ufA83d+j1DQhsm9Sxc2aZXMs0nRxO
LUUxfszX2ViEgBZ2bYK92ecLL29k1s2f8cJsIfft2DoIpfu5THJqpG0NXk11IGjt
QPvBRWCoohvgeTVRFEUZFb1p6oojIZ3SwO8rlmeVA64GYDTBAjnZbbJH/pjhaKKw
52cG7tsY4X89im9SuO/nGgIjc2ECN5XUeuXzgUX+FkrAM+ZxJwFPhpHRCfLECKu4
rgN3uOTiG3WWxBJ5sfjEIj+fVp8Zu1Z49LHVFx5TDsr1ZQqtKGJ6YOy/+odDRTPJ
frF7MPh0r4XSEjUx7GhhAZEOcKJylheeRqANepsteTo/NKAtfQlaxwCcghtBwEPM
rKRB/0luA4/eY7Q38sOopX38ptg9Gw9yCaAC3E3bIMpWdLaeqt+Wn9FERrY/NTWS
5p3RT2IDsYMjRP5nxHsrdL1so/KkGPuWlX3qWRi6XUojC0DYTuVIr1Osr8U7qsDV
UDdHrH9+H5jwwsz+x+EAITTNZwsLYJACD/fM5dFifrTjuYyKBTSbZdi5soYmSyn4
0r/8+RoRnm9XNtSMiIZkESET/T8oRWfdqsSTCukJ2NKAi99wvMFMM7tHFeuCWy8K
sDs8KmkIbf5exH7K80Sz0RADETn4Uv6VqOhTBlA0vEiZZpvu5R2Zofk3YI5dUU5y
670YvJgrTLfUIF/cCw6HkrZS6JEi3BEw4LJO9OP4KcysE2cXUQro9Fc2ErsPS2BA
TqLs+1q5D0+P92vHDIDLxAw2bZFql8KCKCLdMyRxZ8y/fqY1ZIMOI6Vy0wmJ0j8N
ECAc7NR0pdYG/UfwcgTiqyTzgiINW+trXuU2MzOh0J3LHEXC6amfvA/6/Q716N4Q
ay8kKc5Y5NCzHMKwGsPiRhtmljmW/d+ypaUAyVke9Gag1sd9kjSfLTykPo7BMsQn
rbYKcQvSk24ujbJJ8hIs9Yv6VoRhxamGDSn4d2Tcm6bpDmTlw+mvvVWgTPtdMc39
EaO4nEdjZpH9hhq11aG81DhqnQEZLG02zbuHfqWNxnA7+eYYjFdJCtBDD0lKQpfu
kZIDRVNGTbgoAiARd3iGZ7R428aw9/mkg7aqs0YCYhPOawGtsERgHyJZfLQekxTq
hHXxIata4inpur+Idtj7XQ7SUtI1Q61kpEXRdnA0nIccR0wx+Br6gjTaYQWooZt9
DKV5kY/P39CBiqSO1VdGNGbzC0RuDTusdK3D9L0CzJ+0v2xC/1YLXWlCiaS/6+Rm
5sfMQWA6SPQfkaywo0DgUFBaoQ0TZaqZnOW2yRYOF2KIvMAJSOhp8/RdyMBLXX6/
3bQkCf6TS3oxGhGuR9gHeuuNAPf+9tWo8a6FYCUeBfRMq93qx3VUa3t+iRrdqSx4
cNGiqLlzjPfWo3xvcxMcWTGqP6VpFTbO2Zv8sKBR0KKl63QFvi71i6KLukQhV5vy
xOlbZ1AKcNAICZyOSf2ww32+8JB/05Rn5uXkw/Wq92p7A9CMTrIDIzN60WLnNIDL
5Umrv8+EHB4luxSoBGF7xoS+QeKczHM4Z9RjPhJzldYnbgmRUo772JEp7Ao2ASwm
hKos9MD1ch/LY6UlqlvzTnw9YrMISHLCyS/3E6XaPr/gZmZh0B7jyyustom/mhZd
68GF/dqdQRPuZzkP/qEBnLXdegkHGIoIAZ/C3vsJ84pgo6CwCIaK07+qMUbJz1XU
RIt1KG9T4vNAIhuBabY6Sc5rMfeXCr8JBKaC1ziIEc+DysVVfPo7rds4kQMNyzvm
2Ip4vxrqWRVv8ExdXLGRndyLee2VO36v0a98+C/a43zMxOqwHyjo8Vdzw9S0yQqU
57psde4jhl3YEJgFvLOQEs6WPgpvGRmp+c23ZbAomQuN1VmwWogDENfPCVqjVmI4
fOFXZBIqZ+u5YCQs+Lxrv9Lv8DFUGnN4Dwrwuz8D8XyTZYm8kqeLQrJ+E2qsai1T
TJth7tjGNM0Qdi6HOMf/0SSfAngq94pXuGxn7gQ/RT7GchZlM8is5HQOjh9LdY0V
AP/wB3EVZS9Nd4S1chpqvkFFRMJ0qI7c+t+dO7wtfUe12lsWEeD/36BIJ/hawDKB
U4U7bEYOePiAmLS34aar9ti0c3PWHWjmWDt2t7BD/qRfyxF+mL/+CIlLFoXMhv4s
w1C1QOmbBo3odEK9VwotjZlx90jm7z2xSGeLI2yQd7c+DYzQ+ItC6mrBEFthGkDW
k2x5tUroznRRghqwNmVo1t/nZ8K9+Mto0HEGv+7hWSFsCndsvtNe4GcPpgMBR3yH
GIDekrpDkOGTf1hebuaYLxhOPPf73MVGE+2DneYMyOmFkY5aDbfFo3JPau2XwAWp
ZmDrtrbnLn1bulgPbYU+kQK781GlA3B0Vzkmzh5mAHfir8rneMAwkBk59rJTy2uT
nq3sG9biPP8AEHO2o4Mu+eU5SHZzmQDItf+w3byUr9CCiWpPtDPnAUuCrc6YE76q
vevSAdJ5170kHpdzKflc6wuQ7evYrVcCE9tDh4BDOCazr9Na9E4mioCLEN+lgf3O
K0cA6lnld+SuAVTHYx1aonluv6D4ZoDng+5I1EnqlxFMKJjWNWsa/PDaUgSRNaRZ
8z4OcR74PEHXtrFwEDQvZNWFbi294RPHkz2CiPoiPty+Fso6S+MnFYBdu7v8CWX/
BBupToxHjfnVwMLPV5ifO+jHugPE0IQVxQ5QR3NiNwU3m7itmKus/zFj7hbqtSsc
QIZYafJG44TxCGUAQxpTbHNl0A88gGBz3FFv5s43M7EzHenfTt+faNMg5wWbyC2+
h4aAApxAqIlWQhqMdgZ9XvdTOSZspjwclGhEKEtfMe9WG6yM3k2Sg/Wcfb7EBxIP
ATsYh7pKmcPP3z4bMR8Er6cm+accevnTibuFSSioTEzhhAPbcjKsMmCp6We+FQKC
YK5YVWRTofzjCZ6rPYyyNlqIaPERSCHb+pmgLYAFrGRsMdFpHnJD0+qPEgrBGNZM
FGWa6EdVFc/RALCHG/vKGCNxFmZDIHMWujvP4NyAbaHOM/RJq+HuKEnUaOFNtcTO
fkmZk+x5RdnYP0Y511e6XExlbjzjmlVWRJrwWMQPGThSoUY0GBnXs+EBw3F1yU0x
8kei/abXkuIA53h8iO/ZbCvrBGt1FEIZaP0FOK2yROLyzjKXtEg83ijAxDLGhH+6
LEU6G3pmi/pehypZQQjb5fOiGiko5nmru3OFuKNrPeGujnrQ122977wpcouQZwjf
11HE7shVMNl/CXFyUrM9985+5056H4RmTAQowXi4Qgz8sT9qNVI4sd9iWYrj1myK
pZAHjOraSah4wsFWUdxCqhPP4cQfhtOYQSF2HlNymTy4R/VFjKVT09r/JFAdrHu4
COTuweb2cKU0TuDJDo/+OkU4DwFoIk545P+RTPtb3X1MZuFg+X8SldBgGXJ2M+9u
L7Y3JHrB5OhP+U/aTYnpW19H712TLygQzOaRo6vN7V+kwJUjUd+ojmZ8HnPv0B5D
tC6Z/V0NGuWE6S07HNuJio+xtazc0tb63Dv++KtqiOvJtSspvUkFKsCnBcf+mdQC
f5R2HSd15R6CmJdNkD8VpePywq5N/KJydh+BpnUD4IWbjyMlG/nFY4SVaaltsCCP
it7sfu7y8jrvpExHnqKtYi2fWF6yIk5UMMwKIS0vrcqFB4qTaVf86TZhqZfCgPz/
adEUA2qXYQOkjlnduI1TO5qH7KkBFT2F2invK11Icp0uYOnFyEfkV98FrV0s1Svo
TwQjkLaV1zQ4b87bBQoUT4lq55Bp2ffk3Dc2ks3oVFvfvt1pCN0EOZY5xPOesWJM
OPYTGFJpTnSHL+GEVYBFE96h72OYvbPT/CKtMWksUaPZz3odJWly2RMarLMFd8c/
41pC9qN6rQmrN298XPCBv1nxZ6NLShvifpRfasoTkrVR49j9naG1qjGf8A7lXDup
ow2Ir4C/59weW5lzzr/TluyC+zL6+y2Tr4Pr15iq/Ih4JEl/0B9GgiHpDJ9fi1T7
lUZpXsgINP0p1XRYmiJvkWXveZFWic0FHsk8cCfvdvPsAvTGjhfwHDlpD0yMLSZD
q+iF0MO9MhxF6lRiE6iTX3isnYxnG5K6Ybiy356UykJmdKLbMROEi6ioPNeNGfJH
0asjtY3mDv9eKXMvYPXNYTjpVY+U42MnlodVrdhnWAHt7hewN6AuaFw6bKG0atwQ
mOKB1Ofqm+acS3SFoUmVrQUlcNFXptkPKu8dXXs7TiwdaFlWK13dccI5A8f6BCyY
fpqNsSWs6BlISljfbSHigHbQDzzEs7leHM3Bisvgu33mrkAbeeePEOFBsvqlWsmV
HJCuNiyVQqMfRkernwzhrdobsNiBrqWGBN+OMDuXZysj6+/arxEox3DI+2ZHwPTq
4uhh9mA+MDZ90aFLZ+OaSPr54zTXZxptkzxaVlfH7V81HruUKKU4MsX4l9fh7fng
DBXZirdYo3hnHI48E/8/OAz5YKkyHS/R5+ONvXmwBZVlyelLxS4Z+LkUFe/um+tw
3PEpuny9srJG6X+Kfih1bZuYMBNa/bQDl55DruVI6xsiyuB2hAgj/F2+oWzb7VVX
f/1gDjdYRsAfTODtV3sQYKcjm+tSwwabvLJH8OaSB1FLLWhoUSVNYbSNUQKeLmfD
PWInsvN6NrvmJKA7pYvdihdEDufC7sdMdq6iISsmb3k72cm8O7kysMis8syZp4FT
i9/VERZggp48Cn9dRqZ7ya3C1k4FfN3jx6IhroRw1UK1LGhSps/OqxLj+vM3N0RE
gtuYieKaNkfeULmtoldSRuia6k2Hg0uw1nMxk1NKutRVbGq/CSLHZvc3i3fzzIH/
yNpc9coNTK+9VNWJyacPBmJ4aURggCPDCiN/V0a2XSDTs/iOkPHUOSgIznnFcva8
jXOH4e8SydLehbZ5sPAJECscX/OrksyJ868kQ0kv8NyxQJO++KLuLNzFzHNjyruF
Oy2xgWAqaXpD+wweIXJQVR+BAepCzhQ9Ki6DlX/L2FmLJ0uXEI1gyDoXR/c+wWho
1HzHICJqdg9/8OtLI+DYYjlcyQDN97gN+GLH1aG8xyaW7G6ipHiE9cL8p+lffscu
YE9HuKxgtNWduNijrK8K8R2vKojvsg9/JW8PONh+Rf9rZTCbmozNEtC+O5FYrZ/+
99ISesG44Lx9EC/6U+X4nCEGMev0lRp4gQ0afxJ2OK6VBE1/6BrQsFVxUEph6CiJ
gMq/5QbM1gYg4qmvcUJ3ocOXiFd3DAi1Qeb1W9IEjlxvcXfUWomHrQ9U3T5ckm4Q
bCKYxwNXrUJ70U9AMwqovGvJ/4t3infvo97XgVipqlc9TShGJNntb6xAxoICRyji
4/vw1bT5TOFNkdNx70DeQtE5eR7ViQczWDZizD4e+9Waa/o40W8gFrsF4HhpuxDK
qQLhTEynuOIzjaHh0Mgc3AaCf4v9y8m325tMeUud9Usx7E/l/5TXeQX0sZYsJPxN
8YcpBGQNfNt2yHrARB9jiqjZThFOS4hSV9uJudsyREf5y5kfdHUuTJd2G9XAp30+
KE2l0qf6y0pIKPeymchyV885LCuNffUHnjLsmkSwlNJizLaL2DppETL2KVdYuIqJ
GwG6TN4fzR+lYBQPIqaFszOV0k9eZRZsH5iTWh7fWv/M/KGccFHo35CDzsAwXfG8
9rdjlYniZUmo9D6n5hEtLIvX/b2YotvKV2BSwkQBLcIG/HUReaHA47AclV/y0JZM
iy5zFbv1FCzmOXk8QCdXpnwGg2bQMbRLq7HfMNeNkTKXzKeKKznTD3Q4j5kk9kfu
fMAWetlRWesKb8SifFXq2iIj5LhNKUL8yLTG3yj1xQhYoBLZyWK9ltGH9UHzjtla
r9lpQrSyvs7daHxcW+D1XYBDNohQOYJ98UJ8HVx/KE+AiOSqgsYuZKY30TVACPKx
uKmyH/lsXgRyBPSiSWG3K7qZYPW0HmTjOLmeRvB3+OBe3Uahu1C+txxRltqseMtY
ALeUP4IC/Qewor7DNYAi0AIe8ePzndo9683lRCjPYwEKRFHi8jDBWlXd9nFwUzM4
1hG0yXqztj+Hpnag6XqGwk/AK4aVJZz1TkgzkKTWKkCLOCb1qbd4wJwwXVSF6kFl
obCnyxy9fMbeHYWokVNUWOedaKrs8qH2gcSjrqtKMYoAOi1T7PvkYVkbiRb2bxuf
/v84Dhe22ySu4K7Y0qZWTVMB27fZUvxSZlLpQIgTjdgR507Zk0m67LjHE2Ef1Zxc
rZVoYZUoyFf846gN3nHJwiOMb6p1awJw8mKtbvXxk6iW79T+bagXI3iIWi8hz5vb
9C+zCjGIYaMjiLOPbX8wp3l0jYP23pMKONmAeN25V8d6Eq4BkE4cArTrEpK4Zk0w
YJgUN01Re3zOx7ubHFB1aPaBZ+W7NbV/kkox1oFY46zDjzU5V3NGCMxMUz3FKSx8
A38FG2GlUO4nFNspI3/jN/xHPLUy2vv0fPLDuMjDzEO3Drra0rJRuu18iw54lnsr
PgSgLNVBgBuwfnhOwG4CF4DrbnU4QK+cbZW+Y3kolnpulMvytjL2G4TMEmHBXmfZ
almj9jfgOfUPlxjUq53onPiAZDnifuzR0rGm6VvmfGotFhFAoN0K4V4Nwzd2h1ho
jEVRVbD46Hy6cnKoCgpiTZ4ohF1fZqiA/Cxk05ytGu2P8DXdx3iGe+M1Sd6wGtHk
DydLmitpVvDy/TxQaXF4perCdTbnrfbPhW+Sh4HJsxM=
`pragma protect end_protected
