// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hu2J7XGjorVMTPYlqFxUjHvC0Ii4lqGl4Y0zyY1nYhNPeZMU8lCE+517pGWYAg3x
IZ1BS3VlPpwg1Ol3Orbu8KGWmRPFs/Qn82E9TSoK7neH9htMXO1zJuVjD0n6vztV
1pAJItHY1LG1dja77lqhA/FWUnN6CBX/ChM4iE5pqsg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 124048)
qL2tmrPvSnX0nc1ngVTmHR7OaYDG1YiFqI80sm4+JLtLeRbF5TO142W+lSY84TG8
T3PHKszKUHBMNuu5BoQphaNpM+eJkpnaMOmBq91YCX2MdpAUqoIPiVsWmm5YMKt1
RUa5z2x5VzDZjxlBu5HnWK5Kv63b4eSfst8xP09VpVIS/WRSzhRlxPtK/QZTq5gW
lcxKhnuVLDt5fzy8y4LyWs4ALzeJdTAmLvJBg4XrQ/GCaS5KFqRlLSlABhDw1Fw/
Fi1/IFygEi6fsDuI9URauJnX9e/lW6ml1Ns9EtS/TytAUcR62X3c7rnyqZInWfyW
ImAaDTX4AX3SS2bij9Q0JrMVexPF3Bf+61pQS29nQ51DtM0S6Rq4Mew3VRmhMx/J
M0fkrYCHvlHPS/4Cgh7zmyudZIz69rKMzQ7A/KTxvCTX3qTLc/ZfqOt3ILivMVA7
E83hNf5I0/d9a+ESTa+ZaEB1L1QcVJ80BousyGz/eqQueUqEJF7poJA+fu/ZlX+s
8ZuAwz897uEXHJs4gtWUUNGoYtTiCAa50719MlzgAFU+hVcF/Bk++OQItMJqbbSW
ywQt667GGLodxlLeXqU/sAZIY/aNKuKiVdsjCPDgqZ+8x6s5KXH4TROw3qPLcRyM
f2/uIgSOVWSpfLWXofs8M/P1YzAUMc1IfAvrpTFNYVyylpUV518fYzxmV0ku5cW6
mqiscS84vwnfea1girMexVzXoL0e8c4UW6vWMweHa7B/twNGVy+hEOtEsh0tvMML
QJbbwLGQWjioBVgcs77ekL91pPo2aDV0WX82fcFryxvWkUI2cRGf+FWEHrouGZK9
FbZ9KXWZxeBrcKQG2Z1Emnvc28tY2Hdpb3O03FdC7K2V+OzQL4mhd1AqdKFwGqrt
sKlXxV16LoZEaB6xoW11xSYkyGIQbhLnW/uePeF17BpbNcfdEIYxgBet+mBDJgmE
igf/HgWGANKeOJsHqOCdswM4NsZjGCu4EfGN/q9ymFpOh4M1ZnRA851Xj3cI7m/2
ggTnL657hP8+R8W9DOVzNOgr5zlLP36at4KDlaGnVzBNKr/67zIm/VezHy19XvS6
rWupQolaJcs03UkxkJt7fTd8aGO0eWj6IHzItyC33UpDleEAgZDRIafyzP3gyo4z
61YX+JrlMauWiIKMKCR+gZETESAn1zp/ODqHeKYkFRAEJdrc5behGE9gCq3rZlUh
C4GYttqFY8+0Y0i7AIWfL/dQeLjD+nsXGuOVteK/CTkgKojGjvD/CxfFPHyJcY1M
tb8jx4gEOUwugr970j6pLbUvXxm5DGj/+Gy/IY5ZSnTqR+/N/zzTKp1Xw2DxFt/x
T5QOiTlq/0/Onl4HSgY/6oNA/tkysf1tW5F0nj81YE/XdTdQsS+FJKABuStg8ejE
t3ly+oNqfAZfrqXLcSdPfN262OAGJtVzGbXWT6NebTuQwO67uGVLphp4rMS5zN5S
0snaMAWNqHOadtnu1Kwu0hNywHafxT3X/lITWTJDUn49HfrqlSPOWGimuiwpPAJg
0IUW2sreEciACi9Qh1UrqY2KKf2fGnD5+88wPIVXO1xOP4t6ZlHIPevi7/OCnSQY
awmDANIhoM91lF1YXETcxfu/nL46+nXx47m9w20WFFO+iY6eskAAfSfrkn1IPpxZ
rcJDx3gl1QVKzRWLnTyiEdNKt5Jgna1WqOMwFGKV69JV2MsrYjC2LazHbNaK+Gg+
NbaDaV2xVtNm7Hm8WEC96/oYaO73Z/JnEuxePvxZ+M08k4kN5x1RDDesdfInACSE
Dh2U6o2JAyVSy/4WKrgDUV/cahSdlYgJQtHr58kvdlImCKM+2cqCG3I+PwffcNyB
6GmfbmlJT1xDGCs1EkCI/Fru4GjkaCfj++oczLleRoUuXtskKbRxPE1i+/fLHasr
ddQZA2wtY6KWi6jM8JBNGMu87e813kZwUQmXX/sqlrT6Lnpcx6VsxFEYWwZ84ECd
M9phnoS1STvPIH3bEs/53rcd9FIKyd4LUc7x5m00eBfh17DwJs7ZufLM/CiSEm2/
s5YvR3K0pdYOQJ1EFrZv1ztVbwLHuZ6bFTgDXqZed7Hg7HSrDPfEvHhhk6ocSrRz
P/YTXs7VZp7QY1fZvTht6YhZQGJritdaI6ez4lCN5azVMeZVo0ub8/c4b5nJFQKh
Uej5U6i2G27QjZWNhwEGGRoOg9Jt11XV4Oqu9atpieW9OGkfwoKI8Kzm8pjNr7h7
ZvFZO/BlQzZcMz7CsEocQ3pCTaWcmM2V87S64UGTOfO/nPS62cXTbIk9DhoV8Rfr
ggvcaSRNjyivvm/zfZskP2gNrMyb2n0otqRabUyu1B83TensvhkjXN+Xvnx/nMPY
fflC9UBwN5p0/s/m4g8i8o03ueGjS5SoigfnPQHYEPqnKHmGZQ3+FBse1PiEFe8t
m8W3EL6X65bfSoX3zaASiCV0hkFFCM/vn4kFeem0PWQ/gEw5UXj74WvZgw8gWtJi
eK1pdA5Ac30l4aOcDYxObA0whvA6udnKvURMSZ5tI3V4fw/JjRwWXLYMckZSoR27
ov5qctf9lA9jb8Xinkq25B9I2aiRSliGNf9dcwvQ3tFj4vAjKlJeenII/jhJuCC+
7Oq5O2o3pZae+FblyMVcFHp2QoaIorFj/Xn3H0inRpDKDtPgywz3BJzwGpNpcMmp
FYYXK4OLP5emS/x0YWhcozjsqNCNuyBC8F2HvqZZeQ78dpCdG73orfSnphHzs2IU
19YPFbNchiDio4OogpZaDxJqjA6K90G/m9OAmSph/1HHlYWhG0sc1U0K5rmk8giX
ofVNfVfaisBvnDM0Bx2tqrP0z4QqceUKJL4MwsTH5NMG7Ifdq+NC3KHMB74dmORM
ER2ojtQ4hitJZABOIq92icxSiyPxS5o4t6Uk9Z311CLjeADnnIY4vl68FERFj50O
D5fNkN0i0LhMlQiMSKqDIWx/iGBWSDISe7mntzNxQbUyX/UKwDWpsfxa6oS/YwWr
7QxPk5gvWBM64ZXlH8/askZekkvKkrsSLxJZBpr2guUjGYJmf77Uw35vvr/lfYOt
lPm/wnnh6UBGNC7RM/Qetu381OZItF29Ywd46TvcpaKgsnpjtkFxPf/ZHNN6fDMw
qXRoubdjCIQbMpb5eY0fC2B+Gz0NdwVtIPWczqGCVOE4utZqCWKOOyUzQuuL9ZAL
YdD9lqHiw5wAe62DSeU/ZdEzhz7p2+CejHLkzoCiW/13nDhq+QF8MIzbCz3QKE/L
mbPBNC5r6cPPvivs/KCyRka+ONii+mZMRrKnqeBBKCM9BFHWClpz25VigRQ7op3N
R+d8J9HsTAX00n0PvOfS9fb3mQFd9k8T8dMLvACB+BXt0Z33yBGN2fvujKThhQjd
jcjxkjZz/Mt3MHIBuB2lN8rvi7mzQF7XO48IQZVGs4luxOJsudaWtAyUp2Kd00xx
wEbXDO5A/Whl8vdFlISouSq2vpFsddNw4Bz3wCXjcKc86yB7maHZoNgYvF+nlDSw
iV3/GV8ClREj+1xjHm1VhezxafYhF20FEkJPx4nlolygx158z5D6WOJX4uQpxuaq
dCF4YwAQ+/55HAEb2b7ueToig3mTCBqV+Yl18wys/y26AvngyQOKGc3DdSKtoH8W
M2di9BaAqY7g+7/y7QNSxPUYtZv7VdrYtQgnbhXx79bb3fAjRCVWjzrvFdIBRQBE
6tHz9Q56hwRhIegHNpErJENyak0rcWxY3WbpepvFJfYHQN5/GXnwuoh/g7QiMnNe
Zj9CaKeE5hnmXWv4Nbw+BGEb6oHZ/fVnh5gUzdnFwAY7rfVhwRRBMxqa+5Nl8yoa
oiXuZY75d4+/XDXxSY6pxiFOF/+A09DA8SBmiHCY1K20xVMye/RqWvvQswdB8rUp
ZkvpuWGlSZejwf1Bo/dwSuaIKzWzzNcajMsSu+4AIv1qS/MBfswT8qvygnJ8ajFU
rXXLKT7h/0+SVc9/BTAEQAixI+fsJ8ZslwkOFppnGWhforS3bnvcQqFLl9WXQl2C
vnXf3zc8whLvASJuoglbfJobx5Pk2tifPfZABV3NF5eBbJw85t0AHm/rXy6u57Ls
nRjd5htg73/srAdmV1Bs0Gdwu3wrPvKTUqabN1jodsyrbnLlR6ie/OElIRbhCzVq
lGgAhobH9sYHzhHwMLIXm9edkfQ3x8e9vzcZpmOLpSNA2uQi5JgKw4qBHwHYV97E
lTJs0KnqwLa108e+HUo+9KeejPfXlpLrSLsbsWS5q4xrPCh7c6rmILIuHidroeyi
OeuQK1c1+/QUBcewwEAjx11lsMrBCIOQGpemaTPFbKMshUamzO5ZpJKfGRvygAAz
9tcGAjHbE3FWw9mJd2ZycufVllIa7IcDs0io4bUe2WVNTZTVG8GqDDpzQDLdlC3J
GJWp96KaFmlR6aw8OssA2C27EoT6dL16YcxYMzpyKdufM+PxwIEsSrg6Wi6HErWh
qqjTEJ/S5xoPKOZ4cxv72ohJOb3SdBAALUlm9N248ogdJK8wwOuTipSaUk1ky/OL
gIMIieRcbXr4+fEJj2zMs/F4LCViwirMdeI71w8vo+BGq8cuEeYyF8aYJCKQ47Ml
7qTFoEw7E4lUKUjdwJAxwWD3rRog5GPU2WHdMHNDw56LaQpuxiqLmWSMUMAGfFjY
5BNn8zMUZnZF+wFFlRQpQhaY1v+nobhk77OOceZoMMd+fEUebtt2y6B4Os+ZfiYt
7m57BPFLMO0c1Qf637MEs8uq1lgdYprOHomRuu+L5EvpYJ3htgtY/Mf+K2o2luaI
YYaqeFI0WID2XajXtKkQRpybyjF2RnSQHoFffdYkpRgfRCrAogZuh+8bLu9LLCwy
whtLGIWSYyyZz3Ig7FLBNEiShncAhYTftOGsk5Boa9CFS+S7I9uJmZRe0QLVHOZ4
goXx5WOkjcgyb4biSVkWgLM8AJ1lHQKjz6y3UHXuIENCn4dxeM9LTEyVPAJ7LV8I
F2TmQ/pEzhCOdsjWDAm/s2pWgKdZB5kZWq/2etuXkLUzmI1pSk5lXLp42XNrpU/4
Vi9dzwOdDd6a84oUIPWwwjSSK/dl+hOJfcStteNz0Q0s0Cb+U7Y5PenrHnNA0VLT
bwN6S4i10Vj4+qfHFcQIHtAtf2glkZmNuiJJwgerVwZqh6x2qV2GRwkNHiS0/X9b
dEsr6I9R1UgMTl8dxuAqmW0fP6LudmaeXOffze4xdqhhZw/az1APhBD18tXzEbag
tSPcULtIu24hDZktX4uEzdlBrRJjW7SItn7Ybxif+6B8DTLpvZVm96YdFwrveuJS
06TNyVfQVozQ2bZLScb7SAJNlNH/5JB12RYAWV1DX1dIT+m1KaSS9Nl+K4zPEJ8N
hMVY5Oj2G/mVjKlX73c+vBQ6MtxjsiU50Akk66PIj6ury+hyExU1HdjrhQZPq1N7
zZbV2RYiqhiVGvim9f7+yxmGn7jMgc4vFxeD8pUerirg6ndc7knMjasJLZ9IzQ3M
zkaxkwy8sWRSj9JiMnu23K2riB2LoAVzZ+uL1iVhOX21Puc+xhVoMjF35WlhHZlv
7BH2cs/MA+4BuvF+hMo2kolqcAYV2XBmfs4Hb2uDP0jQiy8apviQk7evnmb8NNgw
qOdGMEVVyTwE+GpkaBLMO8s9A/iPUh3g0+4pwMA4U57RIpv7qFafp5qZNrOVbaij
5dTiTEJc4u66303JSjBDRH+IdAjZQ0p6bd2ns6EAJCUUQG9dw+1Jy2cJBU889fuX
MD/PVoWypSkNDjL3cZfEuyNK84Wv13ZiKCAXamrZOxccmHKlyI9CFYBnBavgkUtX
geSzFwo3wEC792yxIhFs3ArJaWLGA0l44R23sm0IZ+2mmTOx/rV3er1CLj1mRDK+
f5T0ZvYV1lEC7LicTK4sn06CzAtgRogFehEfTVlqcY9Dbo/HJIWMErXbz79sSKqj
56j3HRqhEjsQSFCIUmAA/xCAky0q2Y5C3IQq3xt/HVC1RhHBPKQht1RuF8hF2IQU
ZbRDxl/HcTH3CwW0MOeLxM3NcxfLwmlo763KhJfeSo9s6fSM02Xh3nMPm33arblk
zeKNHUJy01kIZxe2//qSPRN5MOOJDprS1/irxRj1cfcn3Ga8cOKssq9Q3zfaKFju
mVBNYwYcCSE15I2rNkHpTPBlhSKtAfYvsFIHp5Qf0Ur6EjAUerkWllSCswYxlFlT
Nvk+RfaaFuW12GM7xbW95VgJgfjbjhY+6gSMMm6RjZL2z8VS5cuFBV2DkN5uA3KT
o8XCtSc7YrF3u5v5dykxA0pFpoS5Ij0UYqUR9V0INhH4o58eJvUFzvauhd4aiy7G
IJ2y3qZt9Qd7wFbZiV/lNHA0NPTTk73dINYWyVJY7RKZM447uLpv3ENAqr6h5/UR
DqujTM+Sp4jVRIWVnDk9/yDdksjQpDLVCzui9Tb7rgiaNi0kI1gCg+AqC3LCJX5U
1nqZxwyQYroLPi3LMQKIqvfoUESf9U+iGa4RLJnZe7Qil3aH7GQ7fgAbL1TTwOBT
elNZ6mRy4GGaAv6KFNjR9czpRAuE02GAUOv6QZ25Hrj5Wk9ZhQEzpdDv7cX7e6Xa
A7ZAnmaiHlym8jx7TF12GGa3BOtmZ4n6XPERdfqdmE6qqhq2GShXrGBFbGhXD0EI
wGR8OIa0GDEx5fCMsI51WWdCvbqpNy75k/YQXqD1n66FobF+JntnIWIL9wb5JNC2
VNldRQUB+yeyNuiz6JXMzDv+/QKFr7/6f8iZMV5dZBCs6b60MTFG+RD+/WbcvTqN
Ym85lNh20n/mlDbrGzmJ1POog3+bYWUTMMaRmthza3S8eGC7fPLErj+tlMO+xoPE
k6XAcmwH7cW5LvXZ/a+Wnq5ZkPgwMiAzbamfL9XpahGyTdibkbuJkbTdN8Oz/3wx
WF3ONFN8fftGOcZowisvxIjOlRPPUI54CZ6r/5lS1/EFr8PbYIiq29TpCE03cOqe
VL8dO/O16o+Pb8NzYzBvmY4h/AJcucoDWyJ2PwDTMYWoGuM4Ps7Gu24zecvNpma5
o9BfW1opHZG9R4xsVRA88WnXIngfMpJqCeHbxvebIWxyecdEOfvntAYBKRm8Kiuf
WWHL2dVwdJ7ZFGiFwd9bgKa9x8QGbbbzEDyveiIfEMfRjnRfHetXlrnzQ1R7xTEQ
NrBp51TiP2K9/Ugrna5axQ9IgdySx4lisIlRMwXYVdho9YWBM5Q+QXhSXSupnYSg
4Ovtn2SqaDrlOVQ7Lp+1WhBZ5YpZRX7xUiZYY6cZQvq+SrBd/0oS6uwE2sNsncCS
WVYGQxsv0MDaqT/CV1KHzuSISwqD0VbpKdlV/+H+Dn8qkuIVtSCDRJpkwZsqz36v
gw66rZk//FpgVJtmEMv2EP1uI8K7WZhAIgIjtYWxLeGzwiz0AwY4ciNbdAAY1BhJ
lP76sw/dcUkizIZhfc1gwdNSFL/IbgQdGRHY+eDNBdXum6qYpItrcVgCxYPqlnlt
fs1Q3662Vs9n9/0fFTWeg0KPA1NggCwIuSeStu9ANfJY4n6jWe55JFB6oEUd1sX4
uRUBwlVs2awnt3Gh0Nv5ZZatwS1V0TRGdORrB8m4FiwJTKkDtVlwdIHdGzx3urtI
rOcOA+ycH1Hed0pJQkVfGOm1xPk2WQHe6/HdByFpQCkOgs2QQUiu3s1RAYCWGFte
iFEnqnyb7l5WnKSm84cpwhkHouuBZgk9yGqcTe8nEBAy4JaO1NKmShgk+mUY2oMH
+XXOPHkNgPAfPUwkQdtIl/xhTiXMmUMuOrDJx14lLrIsWRvGZqDwN5suKcJZZqNZ
/yetU3M8OEfZpenGr9r+SpbgHgp2+jEqxJd/thb63BGCaPytL8BC15Sa7yXn3qSQ
W+opK24b3buQ/mdy+dHozFc5mrcJHZoW/08uMmTH2cUq/IlR2J/9Lentm6H7EXqD
9cqEf47dm6HtIc0MAQ9eUrVHTW4E811mcbzp/aM7Wh4cLsr0nPs+LQqpbdpwQrEn
W3QTuJqoW6oJYgmXeISsDwfzyMEsQt6VC6C4+aoiKIyGeM0UK0upJJqOY55JEaMP
BBqg9w93HoeUZcUoVT8TgpkH6T4dSLNpJN/zLw0YdqYE1AyEkQ88c1nXh4LOhvYf
hhvJczFsmvP1w2xeibrbVf7IHzw+WnYj3Nk2ENKNkYR6ZvMO/FV+1AaedbIXp12V
jpfOGwsI690VCPGHpu8KkqJSKj5Ye10pP2774dSfS9Jd27Xb+nFQYoOVRr74aPuR
iM+MUHzyIDhOqWJBFGGHIMvKaEkIFmCD0EdywLumkCg9ybtPilxULXdm+m5gIUlp
Gyh7tcF9R54ZAW0qD5kWHW/VZZWv4cL7ZTkQvqpgPSb+K09SoFJNEqzmhaDXLqso
gZkmFmaZcdgR9eCGwGYyj3LWP+mpgRUihGJfGYzOcQYhLBOm6vdz8UzKYpmGIe7F
dXCBQSwv0S8tfV888E6UNiOOeyd+hbdozgGt6g9+zNrl9dML2SO0SfBIOyNiCpWi
L6tv0qQFv5RsC/7ibQULJUqWyceOCliK5Fq7E01H7xDyzFzfkUn5sl9OxaMIHumK
BD+KjV+zXxwuK6JJJXu4xkC77bsyhlNUHci5cTEehDH1AsYFSIA+vtuW0oqZa/r4
X+Woi82ZWhbTVmO0E9Xhb8iiZvwgO/nlLRCvPBtr/i2Cl178lJRrBcuCdjb+M8fL
zRkW+zcxyGqEmByXhGeN/2EITcmgJ36M7YMw3DP7+Utml7d+hZG5190r92jQacmB
4fL6Wc1MzpALzOt4EogbxV9caAy4Mxn+iU7oLFz+kP0mwBtcCQ3brXyT28zma5qD
UpysysQTvFCsCCeERyKkGxLK66AAGCuGTkIqKSvSfNVGUJKNz0SnTbLlqhi8TkiV
fskqTQfYNnu6jti9CUMUjQmosXSOgMgdidZZuEF9d2TJOKiM/z3pzGczvEVTeCoO
aCjbb6VwwkmjgCjeErsVJOtbYxRomB68uTiSSGlInKRxDAwsgB7jsVdEqxLOpi59
AUs5Ue2bU1iXdLLWK7ZjLQ4wML9oxFgPrfRP5EVuMYCHNIt7YUASZqUDT2fxfFIR
UygEp3Za1fBbGSrE7h2iADEnw6VNe++FPTsMlcZUnzT2vJxKTghMYO39vg2V0lf6
NSMo8cV4+NQG6CTxyX3ALqdEGSTXnqrJa/jlcGPTBXGgC3iX0IexYCWr4+pqQrpt
psNftK0CsRgX8GqxPnvDhwKgun962Q71Jdppawqhm8RaBMEfzrBRnYqllikX8SK8
n0Mjznl3+E3Jm70eMw0+WuNWiRcVojeojdw/7JiLmM2Y4f9PTAwYUwFKxLpH47uB
ttB2oq6NO8buzPkZkEhj1CCW/tPe/DggR9/NNdLvzxzX9s14jXzYtwNblUQgxUdA
mNVCT7eePoCKGjLx58GuYAYq+NoDk4SeG1jBt/tpMNNyLZrG4ALCv8XaRi2tvpkd
0IOXQ7vtpifocrIPudK2KPeUPEy3YjDSzpawKHOiFMSD5MahRYZF2ybchJqUqFdB
f7p9EPt1JIT3zahn3hJkix6oZOyzKeG4jBM22V6BrRaL3I2/d29gJv5tBiiTIGKn
5RE+gERDbwfkO8vNu7k249Iy41Bn0b+qEjvUV9nWwTX5wqj2Ph6/4EKpzPbaN3IX
mSMpe81J8+OZWNerOAsRx5vBZy64sTxL8TIeDnwfLqN/2yUxiolpUM7A04yLeFoG
0Vp1irQcSOFH6BDFYn2n426uA69eZPp97kWYUOxpGT7A7bIzAwtlZeBOSF/xbehb
l96q28JujJZEnddwkzFkW7FluYHrALmPdG7TMvTVoauhBFzSrOtmvwbJ2GFoD4eT
o8cUu39/AvDQyAc/LaCildE8DT+exgD0GHGJ/0FRIBjIMfT5YbX2RmpqmeKge207
sq5XwKJyZYeksJTnr3gwFSTUORASSmN1z+pcoyvOSjL46FRpR6r0O669p0yO6/6e
FNI7qWWny/R83+IOOoLUqYrm/dLMcjFUKJj4PA9h+qtTh/hhTBULVfZkHToSio4U
YpbQrnWzAjvnG7xDhX+RyIECSAsHS4qVjI55BnWA9sgmFCfzHvZh4hZb9bOBR93H
4nqlm8Fv4LgbYC0yk5hyQ9Gh9b5Uoh385Uo/3ZY7U36JCgSZYFMzsrnnsvntCc2B
GqIoH3vdyIAFKRZm2dPdpBFu8cN2BVwzWc5qUdPWt1AUaosE4j2I5Ha05FoCdL0g
5g/yXj/7kjh4LfbhX9lomYtaB9BnqTZ+TDFt8/tRPcEleCgp8uwg9UnCFlCgVt3/
bHRBNQBGOUWJIobTJSGztb+g8IR04bS9wo6ataXJbFI8PWK/anAunYXImlpbeCO9
VMNTDDoJbrMj5h2vmb3h1vmQnEyU0R4FDCM32PgQPlsNke87KWFu6yaikgzlJp9e
T+w3Lx/KCX1Cb5WXw6I/5U5PNKD1Qd/8Gegoz56CBT0ElxWzu61uhNOrsnGXoy7f
A6CqyuyLJjSLsIy/6G/eFMBX2IRGXRK43xxoX3bNzeXa8qrSOFm4TCwrzgmYzqX0
aX/ImGqLlY8ycxELIZvpkaHBFYPsgC6ykEH0h+SiYg1D6vLmioJl/f40IdDIC1k0
rVJndLZ5DG5Lan2R1kpmGxptESq1qfOLKjdMaOJrO3bPQQukhEu0Sl3eJ9DYDnih
Vj+gLVsaHJQew9Pso4CeRiK9yPEFW+p96zBvcldjk9Bqr4iFkrjCZAP933+y3rVf
gYBypxog2yzQPoSdalcx6He3oaHwdeph7K+iuT0f1tor9pXg3tYOG8a+2WPbUciH
0Lg25gFzcp6r2Vav3Kfv2VxBN1UBoQzADiN8JF432volA89CvkYKaLIRf2DkdPpq
gMCCzHvYA6srJZrdyQp+sFwcO5Ug9iXgxvkTNyRQVDsuso6Qop2TQJeVigA4PQMC
2Bbt1rFpZz65vFHzwDHZMuV5HPDlGwB+IHMEJ98jNozG28xHvWkTQvGqEm8FEXvA
Xi6FxtL9TlUYIGPxSUm4nNUA46qq+FhCr0O1ASr7QnXPQtBAqB5/VSmEclzsPQzb
MswMIXR6CeGS1YyMUZqnDzXgSaWQ9H2iOiqWQ43QdVtVzX2aSeW0wZU1YgITyCHR
ELv3Af3z+Tlt4OB/lFYvWIA4KPlysHWTe89BgJEnmKkK5pVCyFtltiO8+19EgVIB
tMxpW01g1TR3v1MrfWOne81N28VmB2p6vInqO2tCMNjwjjXIL6IXAZXE3m5vVyXz
JJyq8wweHHzZDWw1S96YXG5j5ftr7hz5bUj19fGTsYExgjiywd3iB0qIH71f4Obz
0ICFEY/wcKySy/PMhNl0RbTDf3PBaqgOYZO7TXI2j1lK+daw2dwoW39WgkGUDUHo
Vn0atzpU+/cbq8I+hm2gYELmrNJc7mpeB5oJ3Gwopvra4xmapCqUoBQZzZz626w1
ZJRX7U0sUtF95fAPbH1oNJ9Gy/CN7lsvdzYZGbERCCga5WeEEKd63LLZ8y+jMNVf
cAdTFrXZLFo8mMyz8qMA1F8HSSvXXATZMxF/zzV6LkKKD0WYY9/i7ytIWYn3nuag
d64h5pnPXdeL1GQoRerJbuGsU7FvCEBOlwnkpMkm90Z5V1pdeJ3bB70h+bPNEerJ
FC1AkOmaEe5aww8lF5nm4K2ItQjFToZoCD2yigd5gSC5R8OJ7c2YeCRyZyVQJvRo
/pZYqWyLVrPYA7XHZdvpAzeex9dI7E5uLxn/GJfgi7WtqTPPs48qiGbRIMU5zAP+
Imeg4wgOGZGfLhdqmP2DIQXtRAbzxTyOQa1fokfxM1uG8h+j9xPiCn8mMumhYN/b
Twjv0hFR2Bt5skqxAJShpCdY6XRWdzjgGPqm/OkRveJ/eKbcKsgj4+8l6DT6rDL/
u7ipnQVsD1dAIn1yTptiY84SzpFFv/VwB//qqfNshd/03YzwxB2m8slKk8vElJMo
SxX/EaMs3Du4jRIY5BiKD3ZU2KedtwFXNyDNF5pH1AXdP3A/cbz7xKPtARZTJ5TF
lifuznnyTpxXDtroIjkl2VT920BpWh0I1qXL9N9Kbhz5Zow+9FfuthF/j4IPZM06
vQoDfZLNP4x4NwdwwiWmOvRsSHQwWcTX3QKkKpXqCoC4pgyE7PJzlmRd98disb/2
0gJdMWQTuxx9bjLQ5spn5PlKl5FkOsQuuyOwOZTcmSy0mfc33Ices2RiL2jvWYqt
UIwDAixfMB5c2QVODw9ObBrY4RIQ7iw2SRi7p6NrqQB27nu9iFbE9/G3+lmxSTRA
tnFw7izuQa/V118BaX9yvIll/lmlBnQNyLMhrYnnMkGtRPYlLo+Kq8ERbcYxAIQP
AbNNALaWtyNcgKtTtzAeuGmUSOY8qFclYxu327f60cOyM+S/4Z0/bKgKA+KFE7yq
yIN6I0Gl4YwXxIrZFPdDTD2a8ARLH12oba56RxfYrsH/8+WO3NrB/0Zowlm2HolX
zDMSwOfZt03OODRYr/cGocXlnHOc5VKS7YWNZnz9ZRPcuvmp9cw0piSndEhKc0lx
Rd58LqduVXxBA9W2qZYedJ2NkP4rl8NDntqUxRHqSbVY59MwZ7tmIWjPb0xX83lp
N70EbRVIE46Bex9WZ+e+dtDqQP5YEhxOAM7WQZYFxdM7RNNnZYgbyoeWNYWUVYqW
JrAsDOGgCwXrMpb2thp66M20M26p3TqwSzzMrwCQfUWF6Hpeu0OIld3dw0loTc1F
TOjYwyXCi3p2xfcFFvPXS1K3yVhPPFEDVjc5yp1kjLySG/JRVCi5xfVx/pYqTHA8
8WU3aocRi5Nl6gDcEpzQWURIQlLe8VHKHGbvbxxW68BRLVOxOGTS4O4I7a08M6h4
xMBFRNwpjKhChe8k9N5ECNTCLsIkYba/Xd/I1oJEgb7tdROobg5Nc1COByh2jvUz
9P4AN0JAXdlL+3urtH+ySflKszoq7idwb7NBRnOUqaw+ND0hjCDDwoPfWiHnlNae
1E0b+9amPkzGd42VhnN3PqRffU0U2D3kWe0lD1E033TIpuIUk6Y0S+Y1GQR0oWtA
5Inw32vRyvtWworMFFiyhTd+6f+0L8dPxKGezZ2pGvufGWATTXaStDEZvJZ8OGyw
2/41MZZIcs8J3RM6MXyO3NeA5SlHJIAGpqe3MHYk8YXn86AbuK+sl/fQRYrHsEZO
RJHPl+Mzrss+tWyc4FdHSXm34JMnbKehSN+f9ROLD+Ku3Pb5uguLdlWLRlWA5Fhy
aXVOKNGH0acD2slD+DTBB0Gah1Wxt+KVWIGX/cbYBLcUJXZGKfI4/+DwcASgQ83m
IIWs7YpJ7XYoUbhPmB9Uzr9ugklsmW/ZRFWR1XASDzrE/pdatRIJkwY/bR3N4Dkj
dthCCyZegj/TZ+dU6rgWtUjCX5xch6JRSnfVzez8SflRX/GFSBteAwfzids80bL4
gEVL3W3MqTxXrvyFZArY3bJy8iy6WexGDMJri37MHZk6N5OEN9bgQ6sqJde9aTS/
lDuhXdyZduoKOA2nHwBiYifOjeBFxJDtxcPaF8DH6ER2wjQSPR42U1ec9Rg0itei
ZdCF90i4bwNQWINzqiQY0XxIbQrWY71FbAxM+4ndq5hn7MQLhKx4VE4mPqr3yYjN
3rl07tQfp89LYb2xSFQWrRgy03uvA6J6ZoIg97X1fUBK81CYEvvHeT/hbViQDXsG
6L8Ovkmz5D5+CHYt7EeupcPhygCg6v3yDs/HitgGS9YskJcxB8L1R+RIN7C527+v
EVPe/1AviMU5iEPgB7yxPOxap2ldwQXN1J+RjZzBifHLVDaMAXgt2fvjyx+tqYu/
7gv3WBxtzPnz07XIURPLMEAtb0zJjN3jvHM4Wecrq0VkBdpV/uidZPRrEEiYEc9p
DbhsGptnmWuL3rPMji9OUPzBmgakyfKdZG3LVxD+uDAw9VTzwVRLjM8yzO/uxdgW
QhXrVHwitWzC8be1VvKN5NKZFs8xnNpoE8uHj4Rpi5IsEcdGhf9himsApOyQxbjf
eC5Ckxfk4ei9aDclRvYrHhVyTbDhYDpI++z6b1yIi5u3gQKooIQWcZiIHHzRcvIE
ppliIk3ErdN1VQw2UdMZcJREwAi3nl0G+9oCwzHYDJ1+GCq3Dxj2jLjOarrC1Ku3
g2mIkkpidxjaf1z4T6ykR1iPdz+yEyYqtw8RN/is2xbHGqBXqGcxaqYMqw9FkA0u
bbH2nxijkDo7rpszDnrPyqLoi2dHAzFYWSw+1TMT4LBiRLPypABjP3hUXpgAJvpz
Kktwt3uswzunTrmTlE5V9HyiFSstSgq0dJZapYj2f7hIw5dSgoFJplRCF754WY46
lWUZgWBvqAhXClwr1+cMfgkfAECKBZSiFFOiWA+scho/kDfl4Ig0tPfQaCWTvuad
abWioHwJSTBHedcTvv5H71ZM6PUOgh/bFf6r5ApEFAz/s8ylvrQ+/OxkIq+ezij/
VD65xMbpgZBR5yDitm9tM+Los9DqJ4cfvBUwWLydNzvQt0x/o+es8JRPYLsW9QCV
NUWNRnBr5njVsymlbRnNXrZ0DwBgZgz+J7T3v0mVRpZx6a1gMzwI/3YxCWnkGeJ3
ymYBGEMZ3hMLKQcCLGQWQ1T5xtZ3ZzKilteb+V7thClMNBIHyNiBvONWsE9pB/fH
NadxF9J2QBS1Ls7dvRGtIOJPu7EloDjf4yvmz02ommjL/N5n8+40fXOohkcWjVOD
uPWQFSqteEYBiCahew1LGzAk0d/KBP2Fxkksl0l7mT3cb14LjcbpfVax1yKc63oC
DWJTr1T01BWt8hBJdSLJmoLmrmnX4fRRFx/UvpfVivdFnXUYA6oWf2qgWDLRSHeG
fu0PHqV6x7Wg7cV6BgM9r6WNySHPZ91LYgdjs9QgraV1Hq799phdgRGD3F5fM/nh
EkZ8R/Tko5FNEGhLsTpxBqb/B+8xdQE/58iweHajrqREKiPpW3wwdaPsjfZVrVjn
+Fujk0/+WGZh3vlZdQL0PiEd1smWcXE7NLKFUX2QoTsIw6GI/v54mh1r9KyGBuhy
8o2nS8zXOsRfR35bgQbB1EcHOrZt2ea5BsH3+p9ihSAkj5k7VyJ+qZERa+ZW5TgK
tYwsJPwMma1gktFzKih821gQQeLZujpV56S6MVS6Tj5Uek0R50KMdx25VRnYWMxi
y+0ABymElt5YMfzU/XkJvJwUwnYoAosY+t37/FpulF1IUJzdsIKXGzoJGPJCrpNG
QYasbT0Hfkv1fbEGooWLi+pFseeC1Nz7TlCrzK5oKslhG7iA1PVaHyt2vkmUWiwz
0EEZOBmyzVVtpVllKGvBkGqS4AUMqk8FeXDkWRvtFp9cDOzM6As7I3PPuruRfrfo
OjeDZnDqdN8Yy3CdGl5RfCyskeWr1xdD+KWEcIQAGJfU9yPj2Uyp7fv/iV8JVV9/
Mq3cTH0bTTFED2IyKN4cB/cyGwJNulBlzWiO3CqgyPIJJblV2+yRZ8wWmODfMTwe
nbEzuOkbW2yhVC55j/n4utkw+AIdz+gIhvr/gjxXucUutR+IogTX4pBYuisZ910O
M145BIGk/59gClS7+Phw+YVMPdQL+yd6Qdbluo5FHfyLGcE2tNdulPoj6cEwV75f
D79A3765GS19tgeLlzQIJzbzd2hM7MXYcJ9saJ/pbtwyTPiHZAf/UEnaRsk4BwDN
rAy05lfZRaQQEbMmNxr0ufLPF7+U+P/ewYa4XFrtsbsrfcbFUHrH69MZaA6fT2TH
j7a4C+fp1jDwrbiiGotYszaQMUoPt31dPTQ0RZkID1iQOO0bpq3N4guMLPgqOjHH
JigAwE7uu72Jy4zfSIefmBq011dAOSUR3GCAI1ruOZQbRLc00DWPsuXE+GcK8Vo1
Q2kdjD9aJ0mXacwQwDiH15bEl7DZ2LlrMPYRc5PI6tyKmomf/n6K5mVeVYyaUlbM
5EL45nZJnDYm3mRLohP9uBwEr7EFwd6wC320GILevsFmrZwo2fTy42EQVBoMG8bQ
fzsJ8lKkF/UwzPvmVI/hHbsmPdZXP8prhw56MJQCX8icS+5Ol+N31+YrlL9NJGFR
wejhfZlTDnrtKzpZQdLbM7v3a4i8omEsHNpMlAo1Zgs0sDv1i73p1gpY6w5U3+wY
xc4z4LmN9zP9jI+yvOS9htBAIqFFLwK8Jq9E13WEnWCpJBERENFXqriZxHGjeIwr
8qJn1EpkaaBkKlz1Dd51jIkZXMy1o3lqLTe9fv0MeL8eHzkm/QldFyNxrZ/Pi5Jg
arm2YGyyfuaKtg1cN8WWPqB+iNS214E0ApLisvduENPhOanoLbS/TOfRufhBn5dW
cj2kdjbwNv+O1hBBJL3Bmu1dmnqSDoOZuz9CiF3vdYmrRh03LQ4Uw9T6PHykAI7/
DwHtwvNM5LLLt6GBHMj7vNjekYP3SRGFRXEfwXx6893w3nolJ6YhCXKOhM1m71yW
JvATaiMfqn6kQ49HY5gCt1bMmfj4nolckDPm1Mi3mKS1FEDSp2YZA1bj7cMT1YJ+
11CthPPlShqkhJpW/nkpHlak7Zh14QgeAl0ODun5AJu3WtSllVOimOIbFjCuu4j3
lqpxuCjI882s91Koj8MsUeIptQsIpLEUqR+12BQ+Kr4NTz8Eb+WU1Ghil66YcTJN
LgwW9O+v2F85WKVsxvzUHwLppv8K72qeIBIr5xJ/M9yRXg2uLEFCNewb+rZKbEXm
Vj2zSMuE/EYXrWYs3KFLfcNHpQzODqeCmSQJWQqKsAKSwa/t1250gGWpC0fBhLlm
sIXrNLMsrgZl0IHG/QoEld3/4rJxv9n7C9ZsOgzJEX9+amN4KmNVDhMt9n2WLgtB
2GQZY2TRlPnNz+iFqf3BIJicstCg6vl7AHvCC5RI1t1ffF1R/oIT+tnLuqgs2pTC
4QXZVa7zd+9K4aAeF/UrW/0+iDortQ0WdzRo+vZ19QaUgsUhSF4vswkw/Hd0mRAu
Qi+Xf/rHjA160fvbO3RgPli3g8iFnTgyHS0CdwCORlGwaQHelG47rp2bhmknJao1
ihn9+g2W+Ex79UFZskK2B6sHEx3W7DJvQJTgweaY3xGBx3Mr8Hq3gT8fCUXKJrWX
9S41CeJS8c53G8EqJfACLLEtidV34v+R9QMcTJ6ejHFRBo0WU5PlgND0TnEHcQ+x
VLAubF0rKKAMJ27yF6pqVPFqfcuj+h2rQRxnFH8QCcBfA2MWL+rpo/QMCT/Q/xIv
Q4MLbdJxBNEtC0RT8ch1qcdPOwsIg+oLS9U9Dx7/xyAWSPYLfREugJxuKnjRA+fH
pUXnL9QtwTmWFA78YMqDlrCMjmLm0tNHeOg518wZY6sjhy9wr/NCHWTZ0lAjIh3O
JI6jAGmbFuoCHBqDlG/bUkSKXuLzbmiyvd/74MsWjfxtsrGv92fhqZRRTEXe1BZm
ik74C9CKLn2Ys0Nr4znGl1jw6udmL/7Rx8cufEVgnyc2HF7H58BNcdAdsjVmvz3p
rYkSXSHw/BNhKt1R8KqV6diqBUdhyO1rmafE+Ix6YZgyj0vN/VDT+NtQAXMnRc5C
tZ+Y65h/R2ipS1uJoU0MfscgcNrpTK7A4rfqHEaNTCtH4EAVx0OtlaCSLnke3aUA
TETa3roSx3ZKME+qa7Ux4MF6TJXd97YmoNRlgQhwNkNaN2K6LZOfNgzbIqBSEf0m
/eA9IosgnUjLMOR/V6sG4DHh34ngat8rpKcV+dy9Wo0IRyZf6VGtJx5EBePcm8Ea
nkzENLpufYbX4JTgvw7DlsT6UFUgKm712+v3WfhMiZFwd8T//kP8b+V3uwQDHpb3
yxjxt18kZtHqIWHhfWcaWJ+HPguUccMZjvQ8NTsu45qPd4RxDI3SUJ1ro/Cgkova
cAvsq7wQubbqbWaiNP9If7oqnxixANAtyy9BPVaFuZc3KcOS8m8kCtWOzd3vwotv
fQjp5p82cj/4/+aA6Ajhex/CJLeH+INsNwmOW+AUwIz0s3uDI/T/EMywhJAdHXlG
vtWBptf62PM1o8reBBjT4jCU+RXMBwT75dTP3LKmLUF7vvAa60NsZd09e9SK0wzf
jyqC8xDbTP4v1gXAHss0KO4bu9s7kb6vS90MZOFTI87R3q3LjYlIzF98uOMJqXIn
iBCXETr4Cz0evLXOy7tpKQg85BavKzWSxzeZ0JjEJUDTpKvOk0sPkZkTc7xn51Ng
KeX+iXzL0G+n6yNgaIMnRfBVSzV88ihgS3/FvpPBX8jCVuxgE/TThNIiyHe0V5Kj
gPvd2nG3SHgJlkHCQoTkmN1XioF+IicaWb8EVqL48FhEeByOBlTiu2xSOYJZVuBP
O5uRAbwaSewopnI79DSAiQQ9iz+cWxPtGjCVtTuEhoZ4cmW/o3rhJTyRGsGXAO7E
rs7R/rJyfCI2JJLelBuLsp5qgy3GQim9NmKegeOTwk584cv2xrnQdCEAZfFnCde9
15UuG9w/xJBt5Lh0ruLN9pIQMwKCP8ix1L/LlnU1hoPONLnKwk+dBEirI7BGJhK/
YwVDEFdv1CuzIae6L/Ek9qCR4yC8Kq2a6FxlST4irLDS5tzqqs0hcyiouarp7yir
cwYECK8MXkiuZoLf6vQAUtzHrVPHfSO8wrVjf6CSaBLJEwPI/tyMJKsNY2aFrXzS
rrPmgYwxUdpOH91B4/09jf4iOtHWgbZU7lwx5gUgPMFP7YEaf6CE+ksM6kvLv4WP
bGfqP36LS0X71qEWScepCb3NV7FzeQc4z6iAlTcWXbDMTTP7dZAIshAVXq1shLVw
xnl20pJOk3wZpBnOwP8BOhryXIxEjQC42b35wSe8PS7ws08igA3kAx0QS2GT+FKr
NJYfC7h/tvxsbMv3ohCQMKc6VoGE+jWFqoQclUybSeFgPUfRaN6YDn5a8N50os1K
3U07CE/r4y4krDwxHf+AwhStFsjPowUqnEU9/GH3Z3C8hxhrgSUaLKJAlHG0WfFL
TJcAXHkHIzIf26uwa4IDTEqBq16nDjfHATfk6rk9DAaWB31ViARzWfqGVq0kkJBL
L9dEPz0ujsM7sMRX5zVKLC5Vnz+P3h20c3BDtnB/0hF2HVUfzeRBFzu0hb/r/q7l
PX2AoyBdUU6or3CdqF3bjE0vsAERvJqY2md9GBrjI44N3KbTaoFhOB916ZvKBhNC
BtY2E+PKDHsoXjTlMy9PBaVRModJy7J6mwAxRA8PHW+nVIsXYTw5zvs72QBtx0G2
KHscbeiCva1Htfr0ktyWSETS8XWxyUwo7VsOV4j0+vKlHy82V7dOQbkfoTxIyFkh
w44l9OX0RQvXL/nud2NIoEpaI/VexWywaIGARWP4F5zh5w6jAKcgbUOUQBGOn4lI
RH0QKhp9YIvhxnzX7d5cQhPiYXyFcTAd4jduC947VN8M4+mLuWOsvTFFbxhoyiD1
2uOdPrfpN4PjCNznjY8Bw/SFyGWcC51j68SdtQbp8ODQi2AkRpAD/pmfe/qkwdP3
t2ylB59wNPdbjJZkZfw+3Ppdd0F/Ey1oXuk/ixaQIiBg5HW146ymHChICf3dSx2t
2mOdKL75FmIrgsM/ZPmoEwTohZlCv2y5HqkCj2GBL69VUzLnA0bfc1Lk4NfVKZJp
HG2aREdQWqmPpfvYddSRWN8AyNbPWWmFoxc4aeMxe8gkYX5/i0gRB1RfcD9eq5Oz
n6Pt2BzV50mN++ZZ7GdTbo3qdFR9AOYDUFP7eeYBTNocSx5T0sRaEoCdWHMAmhz3
gKI/H6xvJD3c6HKIruKsBPhbjW5qE8QeU82ihXZoVSUY+D2YIdY8gIVPN4/TXmlM
lZv3XM4LHDJ0dpVAw4WG6y2GfE/FUg9hHda+HLE3EWJjZ8i/oVbeVWqniRExwCvH
ehQ4nQbZn6txlqsCDQdIfJRmp5QMDa5v/frQiWQ3JBcdJs+NHGIwdx40yHA/JXda
2z6gchRkDAlkQoyAuJMkR56rnzGQAKi0hRANkbrj4tjgf5YJdxix2LZl9ZV1LQRz
+kLZSlIVVa5Zx5aH7td787typMmk3suj1zNMIEoQHLVy78rZlK5ss1AFgN992BCD
O2ucWUD/vw8XMLld4md0Fr44mWkY9xfCRzMA1+tDZE4hjLULT/WgcPuNT4SSXMg2
3rsnYikKXB4ESFAPwOtrjNg4pMKrel2cIkMeLHi/Dv5rDvbAYitnDDwioEXGcb//
E5FUwylx9P6Hj2tj07Zu6OUy5NB29XSwAx0TvEppA3OZk3wNUX7yap52PmLdhaWN
ebkzbtr6q6vYw51I3hLOPwHe9IyAMAtClHGf3s0HakCWlRzxcZ6udYR9ChYxEMue
wtrud2abskF5kwRt12YJpfAMHJ8fVPKS5XniXjCivziRuPvTOQ0rlGWZmsZgzjVK
N/IXL4sQX3iCJim3bOrWn1YaW6z/+u9jKeWpdqaL7zVby1aYUuFWNQ3NMYaFy1Xj
2IRh4lagsXGhS8zpWW1dxlZD5XZbKxtuOONIhJXzIS0Tvbr0il+FFxMCPPkoXTql
wxlT28ou3QOWrqao1CnDUg5RuMPCLGm42AtbwXrmbL9pjPlJnxJclGZ/hXSnJTVQ
p5eRhRRM7BLoK5FkbaFrHYzT4Lve7EU1Guarnp9xjRFOk05oi2ITUEGzccQwt21a
6YSCAIGd4EbthzsEI7e5YHDXTHKXKsPojTTuF5XbqzofAk/Vidw2Gpp0DusEWxX0
8fLudpY4wX93S4aoUcaUW0dynxC7jRb06YtyQDIZFhabycRdWjnV6k2SJUaEMykd
1bDlXbpB4yEgtFa35+Xlv9MbsgKuPZHbRfzQgPgChOWcKZSvZ3WZw1BZmJ6lDArw
20K1unFGDBL+be7hKxCrWLJcPHtFvBKTdX2rqCjS54COcc6CG+ugMgeFbt1slRpT
3u24AkOPkGRmiTi4ZMWhJl3rmc39Rs3dapTzGmAD0+AkuivSdA7zyBFm/jzNAafw
bMAOuEObxeAEw6k4dGRUyRUV3avBMfC0TT7WXHU8BmmIUQli7q7MOkATSXuYXUQa
OlXjM+9VwCATW/hC6dAafN0FXXpOhM/lIBkqiHuG3HofdHBhkryMxoaXCQ38ODIy
sjX0FUOA0XSC7xrIDAkC+MxFJiLwExFAy58IT91ps3PYwloNSNBixDhRbZqvl+QH
dXls1lMQWdpkFTZ4Rq18vPwKOi995ELRTxeOAJ/dQzjK1mxtjJkB6KDvlgyILrPs
VTWre2mBpX/uoHXFrJOIbrlyzU1U/0vqdeg0bJgdNvZb9OmouYhdhK+zcMclgmyb
AT+lMc8lcQA/ExTX/esx0bWjjaW7GkKzQ+sqwtnhY7czhIzOF0XpPXm2gusyUryr
2IBBaNN2B4HjTK3Ieic331r/CnYG115j36dpcR3rq02aJ7DXKEpAAMSXXtB/1UwS
qd52xBSHb0slu3xVODbM7vYkX8xeyzVwlpgoT6wIHn0qd15iYL8jz3eIB/7F9UQi
U5Fv9wZuwFbixLmvxcbikDG8gaAsrGy46XKcCqYUm+trgjVJ8VLB0TR7WkA1WAqS
kGbwjwhDT151Xh80noZOIVHpjUFm6LbJaSXtjwV6Tbk8OVaHk45sE7OkquPNQkC7
HJVizvbTOH9YSIRbNhPvphwWHSSU4KpFlnkR9Ll7v/fXZDC3fejx5cJ6HHpxNdY0
mEgOqVyvMIUNt3egbtzaJNWeReFRecsrhVpgMcdrisLCnSGJGYOtqDaugGY+WObM
uFS2rGp7B3JQxzzy7jNT/iA4JFUN9Kw833gexVSrj9uQYqMVpW8FQN9CBZmsZDrk
C99Db44ADF4U0nprGq84Ke3s486tNPPyztxK6f8NIUhrNXbw5C+tY7OxryYGgGV+
KpNQuFEtb8GKAANWeTdTH2AjGtMBoUSKXBz1crP712iY58PScIDfoKKMRtxMr5r4
O/3BnALElbdFk0evt3mxFtbBK8W5WTFE0xuxys/UC+8DPNpQElScwnjVFPCPWTRh
N3RnQ5YPYXk2fbjGsqPwGvcX4dWpjh9FME4a3wBA6EDQdNgkEk3rvtnP8zY0xmGE
5bhDsiYmw/bewvlHCfauDnPf64O826E3cIa7Q11xv4YDPZoVefnAnTMGdjlLRa4w
PV05x4w4PvsOSFoOMHNjZ/1HzOVcWgLcQfShcZYG905lG3WSbjSavP3Sv9l20qZ4
//UEidL0qgK3mQcowNrkYk6vE1K0IJsszckwBg+XD/y5Zhhss6ib2OTeHQYyn4tp
4EkeMRE6TFoLIhF7HedORUTmdcF1FHqxX8lbkX5OjOTdAYOyVruo6I8NcuC0nVPi
M5wQ5fbUoAsN7WS4GQR2DaZOuJ9nUNRgVk/cgSzqV6qDTZrTWlyVMmtGegFL5XBR
dL7ZgAdJW9bI3VSwvwWDR//jdD28dBTtFJts6VIpqxZdUIWkEGrgal52BI2VkQqy
Rim1PrQoHowhlAc9FWTuYfbDykq2XrEZtW8BQTDRo2FxkaH49Tmcde0DyII4pv60
HETQ9lKndsUmrSDkEbVW2Y6ZPXha2WqPwUAspBm5b6KAN7lpkJDmgvMUFrnSISCL
uP5t31p759DeXzY72HLhLOZKbT+vTiH8KObOE8cDKCObpR7rLCEvQnSMAc3Bo6PA
GxBHkjGjqu29ZH+Kez4R8JlzTMoacJXCnsmSLAcvq8zl74u0ot5h/c+NgjkJQ+Zs
CEjLfN1tiAxcup3X6igbFJI8lCv5ftWBo8Y7ya3BAkxtI0mtODCTH0KTo7Le/9gG
iJc+ZwcoXQ1EGPMkrHV7d3tnnkwjuiUpnbPMOr7n/a241fs8WBJY/YRn1paQluvG
tEZGz4xuiWMGFteTQFbZ92RryIjrmpCFiZcAlUlfYFim+F7MS6xONQFjgwvtJquk
XlUmRh2ZQ+0xsHhKbDd3vPe2V+aZ+26ywQZV558MSKFMqCU+hiviJVb8yEivX84i
63fbwVOR+ZITnOsDEM6DJSJ+T5E4RiVl920t3WzPu+7EDACfK6j6hjgMySOEZjhr
ZtC8Da2JQmJx2rFW2DeCYQN8oy0QNJS4MNL8tCEh/+/Bd50M2r1MBWHamXVgUiHS
pM5SNeeqzKOTDKoq74nKeJma/tt+CTl17nIKBgaCg1QrPZR7PFPAYOVMwUslDNS0
idMYs59ELCOESNQM07i3r3mTkQEobUYCGd1kCuB/Tny3dyQbeUygobLOclz9Xw0u
3TsEvbFX9PA62HbFYZgqWJlbiU2kWGgAl8ENWqS6owFaYLRTwqkSaTz8WHf5hyOb
eqwAjaZldS27gt49wCAZXzcIzSlzZnqfObPtdgMeZJ+I7TIUPLLFvmYb6wBsc2T+
rDbf15EAAj+diRx2AALLWXqaXbks+2b2x8yX56lIFSiSa1llRyu0pECf/Y920jMv
Z57azsEHmT5tGVgz2APPbmu02uMU7z79oYrNlH5sETV6xk9jF7buw2+tA7DbrR/X
DkqpA8RIa9uQKHiBvAciwhUQR2ymwqP8VCCMdYV8r2OCjH2pQfAQrgvIlsbxqlVX
+wvvLstqn0HCB2oncZalwmHCoieplAQ54iPihLTbNL14ceixJTs02CALz1vovLgj
w3zXY2cNOluyvzd3I8FsfR3yPmtILx1r2rXDELJP0/2Usrkyb5dtGVT+XRXIkMug
a2LQSMidIrf7W0uip30WD9bb0BaifDffRSvdVLJv28BnJcxB+roUc26sGJu2qlgX
Q/ldFhzh7ZZmB5qKn9y9Il29AfGwEPtEuG9SG+6+nJuup6E37M4L0OH8HGf0df4z
5BrOY46hXxImFNuTK1a1KVoP5RZQznIPT3wGfGX7NMBPJb48AzfQup+Cb5hIVFv9
Y/X43RTyCUwiszdo+LNVgkt9iXC3+N7sfNKdkYNT9sboYW9m0lgZ6c/UCPi4fWHR
xkIPxebuAkiLVl7tu27nJbBxGvZqRS1PPAPYa+fCMbQTO/qwL/IZp9QxE9CMBKQc
rVMVyf8WOqzCKFh4GbM8Wr/Eb+In1FRwaopqD0RNUknOEZP1nfbsBkzTe5rWhmwZ
QBFThwC3PErmX00qodNGEQFKxOoHsmcv3O9GbtP26Vp+O9jSfQgAag9qIXgiJ8Lk
I1eAMA/gk68iVbiNjFIS06oGrG/sqMSlrJ9xgZhXH4PDZVQV5jyO6KC9vY+2S2q0
IBye3nI2zrZKwSgXNapxFWZcRO5LUlhxdcxoxUCuKlZIwqt/AhaGN10IgNwhCfwj
p5zQCfUcqDgb3CEXi2PaOc2/u9hroVKGvka31mJ2Cb1E6pvxk6IC1NDq78u6zFOd
LasGrhOCKA0E3IOP/i5vNUiNBiOxC/ADijLWov9sVEPRq9CL1ja6l9mtBNfW+c/C
t6cR35wu35xNnK91ZcvQYWBrvFTeAeIIlNww0HHz4RKxJdy/9STEkxVfyfKzzRkO
NRnGP5kWScGqBmcSKewfDWMGvDmNFjK6JbwfEL7vVH2BZLVDdj+HwuNGp0UGrB+T
t+OFrxKutz16TKmuj3yjo1Wx2Btkk7xwkHlfZIWQCDeHahzikP59kwg3nIxFXiNZ
hScM5Z+h073qXV8GGWywgSJiobM91owCQsqBpt2SnUDIDOtUmQCwuYm7V6/9EF5A
M9cRKfTADegJJe9oxy9pABgD6uf8qPN1Zmiyvz6pgqIaOYWZn9QBwTEFDpMukfmD
XMW0o9/7b4QdxbtkMV5ukathaDkcFQRVVU0TN5QZ9TJtrEia1lDLHqvI2dUtmB6Z
Qt4zjC5HHflHwI1LT6AO64eSAo8eqaan6AJtQA4hUoRlZ+pc9uZN5CWmpWezcstF
iIOl9pJJC8zjGOw62b7P0Mi1ZUoZmDl47Lo09nMZLNEWbIdndxgk9HQia7WBxG2m
M1MctcO2m5UXL144Ch5Oqz5QUuXEkc2ats/H1Z4o3o4CXr7ikji4N8hnB7Qb6cbq
d5rQCPFVPTN6HfW25OMlftyLy9XFGcd0OwzvhoqMB2rT18UF+rifTm9n0NO+ferV
5HQljEP9xkk07l/38sZf5kZaKFNbLAmE/Faxib0NlR+aPvzz+xE10sWM/piXcGxr
FT1f8lGIMwMfmTJ7P0bbMbWH1js0WUn4eHJMOOOmmysKFvSB3LUEJ37MmZTAILbS
TgEERalLKwkvLIke6DAZU3vnq8nnKDkiNqM0TniMTG9x38Wm3fPFAm4zQfKEQ2uX
IbyUpNQzfZ7AULWXn0Mq7nNC7+OAymBDMM7Ehn5CA/Nl1hJCz4dOaGQefGFUu7la
4mmxmPT3fx/fxZbb3DqzzRy9M+saC/0DOKdABrynNMmwypsLWtNPM12MOm08VkWT
4Vw7IO/GQPHP91y0KHFomrntMqSW9hqgKcnlTkDpWLmf6gfpvmK9AFN7CIgyIClu
Mgwx8abIRS/Q6wXvRSwSuCwxg7oUyIUmMCmYEmWBOP62t3BqzEWDv0p7BSVXKNc1
XR929TErn/D1LoTUNdVpa6yexRJzy/S775TZCsoOaW8wFAzHnp1OhMcGewS0idc/
G1vVboah0tdDu7hyw7ssZOK/lU8AcednUp+0P6Dj76lnrmlZmygXUJ7yzFn+2TO9
IknRp4Rm6lHt0gfaPXmE2CsPdm2PCjO+6WZZDHt/6RXRnQWlwhUH6B7BWr1bcknW
fqR0j+sPR9hrH2O9GyxvPOqeoS6kBizkD4MwEa8TJrgvpzoEyrvJaUz+3xBjIfjP
fzhGyrgCS4dMTn53Bzi+UdLSCKQcR4Qen2XvWv/hJUqBx7WzXYvUR09G/59BB9/q
xbRY9VZWLhn46YPRWnlvKXijlnmaczs8O1vLdlwhdM9uN8gG1wDjPaedkfunTCBa
cQhmgidE3tQFtofkWW9xwMCfylW7Di9jIwjub5+R0VbqL1hszFFyBN5wf6lv6ANJ
eVoYWgC0kDnB1WOzsvXAyr8t+sr6FjsmnW1Q1B2Y/xF+Je8Dv1eootRJy4m0TfBN
wCZDZBFBaCKm8DccxaxCu4oNji6QBy/kW4C/eqOrLNPkx5tMDdq/KFzAGldTJZcD
l0ck5NX+Xfqt63oGzELYPlafBeQKHyC9nzsNuNP31xwmla5d1eE104B1Apw1PhaK
Tjw81ofIZvN13R/Ce+/GlHpLoxdj8pO6nob7iNtWIi1ylxzev2NxDV2Mzt6dsQec
LL4xMjAY3BwpsAXgCF5Da445Wtww4pI2N+h5YxjWaDn0/TZFq6tolP73NF2fNQ+l
nJtPlkCF7n8zcTyHn7y8lejJscEDG8vFQTAjCMT5aT6RoeCU8Izcn1yWyHzJHupk
XiOzDu8YBFEvvHctOxSDr1niuV07Gfyfep7H7ClS/YO5mTgmjPffTPf2F3Bpxhdx
vVgxNgUDD6np6n/UPQgZgP3mDiw80XOQfG3FhJg7wsZsmAogX4N4AEncw9Io//fe
DyTn8vGwefHTKqBR9XY/U5YrqRlUglhXxExVtk9nQUBpyt2RJN7O34KvIJnqYIUu
uWgPEi+r8iZ64N2owjIhOW24JqZnw0q8+W2081X5g+bgL0faVEW2nAb9SZgTcxLZ
nLMrF++MGUT5yyIRDtK0MohvpsnC6VksMa7rf03x34L4rTjhCP/h0EsdIQZvefhu
2y6Mad+/Z0xFW3T7V90IM7TkbtXycoLnVF9J2DIRITrmI7r+PpEHRPUmzQ6DUOpZ
V1t7ip6ePJ04ldYT6zZ4PIpEJRpdig5IZ9xtFtdXcYcHsX280h+kyC3u4Iu4yjER
nHA0db4iMzQ6sjwDcM9sCXDlKaVOUaY8pweZspvAzgnGQGe3vZkJFC0WusKPJIkU
5+Tf7fD6p/6+9a8A1yVTrjKqT6jIKFWYb1a45iM7zl7PSmmZ1jOw8hSs71foJen9
LodkVj6a/QaCfZ6vh3GRk+ZHtv9B3vA89gcm/ETKcnJfmigBUjD11EiOHs4di0Eo
WfX6MPE/WJJKagsG693msT1bQ2QgRAruqXhz+4Sy26BaweuehiSNtqk0NH4KKYRx
XpBKhdAM6F9M2JDN/Riix47YPkKXQDJUIDZZPrZmcAcVsouMrthWrXmuX9gKQOzc
TrrrrwVuO+TdwmH0/ZxSfVUTiv0BRTuLRMQ/uN9Z+hact9NVNqCazzFEzUVWDQXk
pd0LFiGzy+A1nuwxbTZfKNZr0JHclvbO6wfYAbinO3OtExBXCBSlQ385FNzTe5pB
UhKa0EQT43Q1bBCOPrcV0Duvswa/PxMf9OvLHd5pk/Y6iBcnYlMyUkgdW4TEuOVz
jgNsZapD03bIJL+N5ZjjCCep3UbarfLv1DiKsf6bGbLrdMWOyZVE3qBDO6ziHa5z
5bB3wCJbmU9CMrQfo/ssZWf7+72CS6Y08vrUsJpkKXjSMLyr5GuwtAk2Huxz5eXv
lmVO3v+MhGCw5GNBFLF29Ve7uWKL3Z6rpdPByqba6tRSTbPqnC78Let9Ya3ordUT
z1zhZCL0tWNQo3pPjo3QvTaayKNSyFPBaM5oQaUjVWPVec72hHamrKon6Dvb68vr
4M/sEByTTlL3WPtdkJ7WYLF5GmEK6EBj+moJ3ugc7+BMQ3lwhgQFoDEHN9tDwSTC
32um2k1pDyPKupR910D8HB0QA3bvzRK1mxLAveInKGt7leF1rNLb212NnuzoP35a
H16sEFSau66vMOF+XhQJUnUvZiBTK2L9/nzYZAbJ0Ez3kwxmUQ8uGYCABhwp1FIc
wgMlgrD+oYkBF9SueafoKQ72ZLTzWLXt0Q8PrC8llzjFXZ2wNJpPDNziz/T1PrdD
aa1kyQEtpEagm+v+ojE7N0ecfxwNPU3FdpvCLMJhnt6HIME+CSMWYktvpianMN+1
2/fj8Nc2VaMfqBJmQWJHLRdmspOHpoM/HMSGsBPuKpZPrsrc1sQ1Toxu6y9ndiu5
DBIEunzX16GG51mWxfuYewxUM9X0Bc0v4BQt08IG1RK3SAyHaGxjeUXbVPwJJwwV
v39tKZ5GC651j+FqPim573I7nk4rYttfyPNpfoBrykiq4VJX1FhwsF0GWn12pq6f
WenBLrn8j9V792ffuInAXWu+aX5Yab8dZUpg/r6NAHOl5+5MoKy5sPrVZm23AoZu
gRq2WbFGkTUW84mMkQdKOy2aOB8RzSPNGH4tL/NUFo0A6z9rRGnZBsZSybJQIrQM
bBGZ1OMEO8N4B09GfSyoI7Pc8q+DKvKIKRPEfmNq79Gc+77ANmNm6gVh87fmRAZK
53Ur2vi4psOAc8xdl7MHiv7fJdwumrP7Zo0WBkIp3HWgnZA+oXKZeejFQYenC7K2
5jsVH9mNN/mWhIN36pTRn/FZYQtyglL0s8a+VXoHkavLEej/giWMsdjcWt8I7rvC
irqsrcA1ii5YShrXwPjhmWasJRYKNaPl7F8lJCkEOmyB8MnxOWIApUM6lDmI8tvK
qwPTbmnqmwkrF8gffaTriULIpTRQyP/8RV9O7DYQEsy5mBi7j0J+WTYd4vsnt9FJ
TspVRumBovTs+VJvnsc34Qlrb1bX/buie6JRQ5FWPvM9Yjk7KfUAFjxL9h8nnNn2
AtQN5dY6YRhTkcEGHOyVw+Q4jwoYtwq1qMzFG5Q8S94YkUFNthLBuq0BGAFzMWWz
NAk1lWSlOd0Ju/Af3oW7CbrXc9UAn9B1ewbxPJc5HMegUpbVjB8+QNiJ9RU9632f
8THiDd+oO7hLtS3fgaIsUdDYHjJ+A46/8PbGJ349uKykpgRZtSrpUmswIBVNjJYI
ICSApggpbX2XdZK0xOhnKL+8+BBNqkfgzEkuY2OpwTdUTbv3NAvqqZjC6SGkjkYN
CuEthAlQQX00r1k26TLAWGvp6dtN9Dot49f0HoNlkoEZLte8OZ1JLt4ibSkrIBsc
8A+PJqJCt2JY+TQc5sRnVe9hsX6XJhh1R6j/3xUCG3vTq7a4G08miY2Vxw9rh3Z9
BMOrxrFT1GuLfD3/sx21vlbOkIGepBq0p58J0u3L2dzbWm882GCEI8RjjQRnuA+L
n9DziNK8p3stKkDqKKHqNEtzUwk8Bh22oPnk4uRyTLoXO2npmcqr4g51sBRNE+x/
EP3jp8hr7WIvcWnY39Fdwz8LvQEQX6l2q96jpyVlTDwk6fTKgV+95iAG4u12VZJ0
epS4Upw8Rgvp+kjSMzsdFUztDI2vV1BDM8T/Ca4AK3SDs27ViZSJsl0TEu8W0nh3
WYhO26j+QlbJw0QFFagUQQE6OL20gto4jQcGJWFHFGAvEp5mZ8O4CcDqmlowPZ4i
092Xa83LfiVx+QFyRxYrpHgMagGjHQWzU9+C//579VyvGzTIQxk6r3HcizPPaWdy
NHZhtb1U1ui5rDyuZaKYjpbdpLJlMxwjwHpIDQJOFvMw1+4B7wld+IiH+Zbfffrt
6wG6+jGAMZffGr1YMgi/upY6JT+JfAapddus33ENH3KbJ5pGRGADB5Ya5sGU3w6P
83Z4XkkvLy4tECIDqz5Qk8AlSbpL1nCDOJwhdlakX+9H5GVxwtxiMW8Nyx5s2Wzb
G0IgfV4Jrld4O55CScJapfMylxA55vqhPRjNm3TZXZaB+Hajm9WSNX8Mf5r5WpYP
HQyL23pmbP3j4PrdcqzPGLE/sZ5BQ6hjCf2INq2kkSjUok6Bsjw2zbT0ElqAmNj/
umUIw4KNbdbyHryQ0rMLnHB7NeEE+jF+JfjAtFWKi1ZUbdpri9S3h6GXZI0XKjt7
b363ExEt5JHSPFdnKj+IUQkyEshnJ98A9lmM60RcMVZmzWjQ9SFNm+AbB/lEjTyc
FHcwgdw6uV0J331Wxblh9z0nmCLow9DKbaco+ijQYTWsUC/i3TUe5Lvav+MWSb2d
rlhGrpeWmbzfnJfrQ54qWmbZ1bbpoJmwm0438ojF90CCwlM0frqPpwCs/eF4DhL0
CM+xHgfpy3JYvUnZtFqt4aEs4IWmROTyeOKxFEYnuUR1KnlG4TxEyJxNDfaYulpg
CN3PpTuwamYC7mbksD77rfTuJliQiMrSwHnjNDZyfeiUCcSHXY+urx8aITmevdQe
dttNxvC70FesfPVMxVllqb7LG4s8XhtKKEtOsjkUCZxWLzdXnhm7TjPwQvI9biWr
qM5KHcQnHBjkYSD+CZRodB1grRHXW/UPO4WJp1KA+d/2/Fv9xEYQAE7/yjTfy7MW
yNvoVcDfcGK5zj7ot6Kiyu72Q36ZAp2FzKEb1zUHqOvuC0C88p9Oz303n6yr/haF
3Lz3anW9VHhbbhThEXah2eEzzwG9dfkyxeFJQPxiAlo540YqMsPFgRFOCEL+DL3v
S9/GieLtaFVZsDzr4TJwOGf7YXH3OAGw4N+t+eSsGEwIkZc7AZVoCeBIDzN39jQz
ywizEuxZCAKCT8w6xJaCQoeC2iHmzb/8wvTzLHvl5wx+Rw5DZLE+mYkrLxuWlygQ
yfRVPF6y67hO7p465dANh07ocxkk7r7VFrMYPoh7NDY+fLwR7APebJz0HrqpZeGM
2xdyAbBd8rE5yxYSeGNgoIw9qCLppxfcyNZMLify8APf95A6h7PYcMYK/3qp7jT2
uHqcQ4UAGePGFNEbu2bPUV+yF2kGw/6ffGL0uCUZNkzHvEbNOLsGa5GCfde6YEZT
zsHn1cWBydH/YyxHJzPk+fUsuZ/wo16icUmHp+/qQiPoAyDmIkdAjOTGXswuVcR/
AXUe68eGhTWyU3U+Y8mMGmBOhu8lU32Y06mDJSGjVJlOytsPTFA7H+MCwLhu+WTz
EX4Rk0kCvkJ+jqTZezA0sWsTuE8gAHiu12Pf3r5AQGYvDZ1c+/wNQ/fkmNXd4Kgc
gEEQghGFD5h+AoSqB2s8PAohb8YvTKsTCqzIQMTCvByYMJGrkQ+o5aAFQbv10Llp
avhGa3RJoEA8chmTQ0ymwteBGc8h5GiQApBhCQ+vDdctfekT2spHaNSP9arlBwd/
i1ZxsCNxdQa+dshotXIKGmZpHFbWlaAp7beeZ5TQ1quDYswpYH1Jy76F4G1HJQl6
LEI88X+damDK4jy8CIsEY06QjYgoteBGnAAYspFORs/O2AMbTUeE/X1jMdd7sU/+
oVIlbzh9eMAEt+b1PBQ/wiBi8O49kqvBbvCF2raQdeFPAtnFXTbTF2wcbo61fuLq
S9njPyIW+6ird/fnenQlZfIE3Wrd/hN+CYJxuSfQ5dnStubh0UkCB4ypDAOP2S4R
E2Ako1roIOdDD7OWihwB+L9s2G3dRclwvCJVoT5qVQNEfVytAxC9JFwLLT4pNQPS
sV4ZN1i6P5Lj7wzHHwM6rB6VP8PUZpqirlWNpYAF4Y/HvDhMl2E/U9rhEHlRf2fE
+c21zF2RGuikfTYzI9miWPNinBk8QDbFMLmNNMUKqqtZB4FQ55CV7i/goBFe6QIi
mkwutcM5sHOZfoewbUA3aaPFg1VigxKvjfqNtEHPn1MrgJa2B3fv7Q7q/RRy4P8E
gx/kgrzyoaANGZw/5WlxEfeko/2WOeIf9aHeBi2Qo9GKtRZ/VaMaDTbFPav5iQrM
f/cjcTpd9kVGFQ8yjECR1gSLo9b2x50O9pUGJMmdAhPl6xoKbhX8ZzMbYkaSsT/2
yP6m4B8G2Em2dXhyzTpHRKikGuW9wkX344pBxdfxoJLw9jP+R7lKqXUZEONQAlz0
qGy87eflGt699OoB7D935E1qqt1p9iyhs3tL87CmLRe5QsgrXSlPbw/B4IeM8nRG
o3tvjt0OKX88pOWWRG72Gx3XBPoxbNOlpqdbdcp+i31Bhl44Sjq5JjPgQS25i9W6
vdP9P+o81DSEdAcPqN8AbjH4bbD8gMir66VVakRSDlM4dOL9QL7oCriziWZTFnud
Ryf3s8NpRx1IC6T1c/bP8VHtGEH46bZlsAnGxnWnNDUBafnsEJAZhPYL+r1E/119
hRpckPBgIH2RNfkbRw2Uy0dsATq+U3qCXxV/1zrvsnr5Z4e+/PDjRJjkhQN3m2zp
56C3P53iWKqVSAXWeJMUALPi+8cIEekXp9Q0GohKip5jy+xbDYxknIaOtCwmYZNa
rdmFvlbAVUM3MrLfnrjcdV/rROl6iMGc/Weabs+0+kZxdVEro93/43Vd8qjMUXls
1sfoAXjf8RIQ2L6bFqXR8YFDj0LRLFobrn0SEonEk/UHJsYB0r7HN72Ln/wXJdvY
VeBBJafzKrwgNXqnAsPuAZmi+8wjndS7uXyXnuu4zjqo9r8zlQh7tAegr0o2a6bN
10IvGF155c+KoD0nDjp4/UYm97LmOSEV02zDYwIif8IrGjFYvseMrlbVpfI1zMHb
GeyOT1qZ7u8ryEjGusuWJU5r/NMh5O1N/GE47VXjSl6AVdMkWn5cAN2E298FiVQJ
9XpnGhmmX8Vg/5sSgJ7ZFBMNu5BsS5jZkBy1Kosc9VtrqXPP4JgMJIFXKumZjHrl
dlzfzWQaAA+UgEJt6guWtk9RX0EabuIkY1jXrF1kYyMiFuI3dpTyCpw6uOAeiM0t
3RuweYuz22eLjmAtLXjGttggjw0nnU+BUiOKG5QtOdV0PS2fMo7LWA99OkpomJn5
3PYDGlbMlgjyZwRd7OcM/YzYLic9SxI3EBWqYsOnPB8eelBnmRUahk+e8wbq+FCK
VUs8a2cWrfaSM/4VgYCaOBihgYaS6CyCIn5dqPgUNGERHjVhFuOEhmv+yDkC/WpI
TlRDtfpVNKQNSmnoYaZI9wC0d0l/9zDa0xGHkehGf+uVFmZirftomO6bV61IFvk+
wRNr3Lk3Jx1mrJY4RivumrUtjW9jtshhMEmPTzsobF9nrQLYeEhOsqRnX3Z1wLeU
EmVvgQswBs6nezlLWrUlqxtIZhmZJ5Kse2pIVYy7MfcMYPyDKmhmc04S4IZZokiw
AwB+PaYcTdbnj8l40DPI+Qeho+yw+Ct5ByYpFRkHK+xr0C60CEzwjFCZaUKnhGBQ
Y2ALHBjodHL6sTxC/2buntct/EQ7z+ow8mimrRjrKQ0tgTxQ9DfzciaMHVyU0U6i
VAeI+4rInJmZq9f5iAnPfaZXSJLFiNHcQYVFju8wgcsrfl7XF1jn6TFMWwoKAauZ
eqUNFOhgkAw/didtjKzgZ8aGopy4gPUZZjGAo7tyi2PDRtuUEojyce3/EzrWDyUS
6YuJo/LQS2tddCBEH8tevYuqilVowgO799NcxZjTs7FoszRapZwbBeV06ln/8h+g
mNa6sbBIqUC8DFcThZX4p6BEnOY6Eia3hYuYZvfg621r9agEq5UjVTh24zqIkAZV
w+jug/2JSVm3+uMUg8D4F+xEiJdtOFX9nUmK2k594dAalE9r79NsXgB0TTStVVUp
pkm7EnLXE626VVvRLGJRxh/KdTHmufd6xuxGLgA+LiEUxK7JDOZV+TfLIJmjZk1S
V/SKk3W0DgnB1ZEKKnW22wQgkxqvaTZvWd7cjZjLuJHghSYXXfpc0b4nfCVwxwUe
afJvzLjn4y7nMWiNp+zcf5e62MmobnJVkQmdAsCqT+klo+CGu4PlHUZLZR4nKM7q
W3lSiyhNOQR47Wx83oZyLZa88CYwxLrgcFjflHjiwap1jnQVeOvQlLdJQHsd0Swc
mK4jXOsmju5YgGSusZVJjVDrWM6/y2uaWyDJfvxg72Ux5NpfUTVIVO0E7RJlt3G1
w3XuFWSHnntNGJcAlFNqXhVb9kAxFoJZq/JuAMn+E9EBdNMTNwh8WuZbrxIM93gu
hzo/9q0XP/AuKgzzSWNY6zUPpNhYjFdN/FhG1c4yIlbd0cuZn0FgozrKiBDFYim1
54HF9YjoisfvrpglU43yWHWlux1AGUrphhd7LVRAgc5tPIgPK2Ed0pikRV54KAxg
ls28Mk43TNMZAvpMl5c/rQeHH9QnHI6q15lttyhCyhve67AW8fLVt7RPv3NF5fLx
evncBWm53sJU2bCC3NIUEKHJOxTECbutZSatz4hIFAZYZ7b7frdDjd1+7wZ/RmZo
Wg591IXJ5gn95eHDYrLyN7CjKdkT3sxO8sqyWyxFLhglfBrwzebycY/8XQ+4fB8k
7aPNkntm12E/MBLQuqPNiolkadbR0VTGwsCK+tE34zPLkwC6r7qnwOkVXuhOFeIj
LKE06vnk9CqjKsAhBdNz9NH4sOqXEQ9aavcOsVnIMSeC1K+csbDBLgnhcyN2gtfK
njJDjNGL2IlA7ExfZGeWkoVUhQYjRJ3lNyV8fohnkj+c97Qu1A/i6TEESYlBWrjB
+5X2pAfYBFgOS+Z2HeylZlnfc+wE2gYsVFEwcIYjwy7mq/kUDqa0ddW/lo2zbZsr
JTEPhsghfaB4NVQKgRWLavhgPm7lCSllu/icjXLx4UVTbcR9LlDC540TRAO4Gp3M
3dBHscbfyVhSrRfjPb76hC14m60ULeZGC8txyvxUbVSXgqFiiLZ5uOdCUMYr6dIH
JiRRI+eKxhLPYDzQ4c75tf2ggXGfAxFZVNuoXCMcv1ZoK+6Ue829yXraLjqGju4S
+Oj0bUbKR+mqz+gThM8Soxv995+6clbGWMjqNPlRYpz/dFh2wHTJqpuUnmn2p/Qc
a1L5F4/9quPYJ+Z1GbjJpWZ3geGpMKCCrG9JrvNNrvlQtf0Bpn4Mgi75P+IzAlGi
vibptf6UgxE679fhToKbMgMvYVzr6SWbKbm6tKHD81s6BECMe6oG/i1S7XNpAuxB
QttrTCWXinqaiMWQ7ggp3d+DbgCcRczhUHI2flOcCCukYwA3cKFc2VfCQ47ywtC9
8e2HBAVf/iZ8ttpCc2ulUnzL6FY3cMt1GTajkpc+JYR9wVSKxhFAYKa49G5Tsadh
bv4CcOajuLhi3pR8PmzyyHRuVQuqsV0EtK3tABD+VQL6Or1kXUPdH0+IS1tVQQzt
dsMYe1Z5MOwfLOOnijHCbSqvffrcZqp1RS2RIqjnwyXz9Jp1v+hxF8r1f7118o02
sI9x58foGGwnWqjwh08MBVDnvDsXdhA/lwDBNpK9sHaIx1WeXENylNF+07kGuD6i
/FyPfcWbAxpcRzziI+TdIu5Ysp57DdoDMjZxPaKfUMPenxAvxCAfEmNRsJ6oLAhv
CVvoI8WOxR2M4BhItBavgeLFpu+cCHYaOvUTClzQiRJAbRy/SILc08B6+X9iHkbb
66LsNl3jDruI4orsfK0EZAWzr3I/0ZfdIzGg7u+dViYazMAFY4AR3tuy8KOGOkrY
yQs/5pUeqr2BZ5mmNK/IVL/sglL2XJPz01lTK1t0hwMsjMmFNHQlvBT03Bem2T++
93kyqi2hkhVKHJ1BlqNG07fpefPt6K3UF/VcFyQ4TAoleFSCSOvxKC8KbdA32GT7
JCNx1kgStI+f6FGeXSCZBv8iPQhMk9tI6vSTmrla8S/sx33KEz+XF5ev7CLimXhv
BjxRucEO8ZHiuZm37x6TMTIm5Qtq4VPY77vbr0OPSXO6sVDw5MUkQfMtXGz+L1ly
JfbDo/fEd1fAaMsGESOPquNKTNWL1HV4kfDQ3OwgbGTzjf35nLaPQM4eolnC7bAS
mIxsjo8eexg08DYfgum30rjVcTvBuGD5UbF9uoOAogx0Yjm2JunfdVGrHrSmx63r
87BOJF9oDZmB0pAidwTXgafNPzg7kOQ9iFuY5MpQ3IaifDU5xL83T7b75GPHNQoc
9ds+SrBwKMjtCkUkBdd8tmEA/OTzIUJIhyJSrVZcsvIHJLCynkOLpihhJfN0u90o
9dtE/eYysiAkB9KXYiof8cThg7dR5Sm4k3fu2mlP2whOd/hFWdZirU4ClHib7COH
K++lGe5M2rfDxDPTyHprazSdeJNmkUGruoXjk69fQadyhGGdG+FqBykptmUhB5/9
bH/nIqkWw32HUaODDuwIqAOSe3o6IAzoWXgpyOrLYJ8gqVGKsfci6lkiHsDQ9u50
twVxJ5VzwmOSnS+PftwSwgqgXSjlPG1MYteBBCy+BRfbGBZuQHbj1sP94EACsT06
cWsc/aNjvTMae7fWjEOuOiKI4t9LZ9qdJoOvRRRoDzbIF7xYTWfV2XkYU4akcgDa
OTrAyQ14Rp/h7I5J6FAwMSl7xpxieaDzV5Jz/nJyDTaKHGUVUZI/MIvoIKyz3H03
SfTf3imDYgR4pI/JGMUyD1hUj/4GX16cVRzfGZ/jPgRJKxjYWl9pyQ9mt9omZoJq
0JToja3sYac/UCLq5riDuiGmE/PhdqabcgnHzWUtHsA1pDQ6UrXA5DwFjzXcTjJz
UOfOTwnpyBN3FLHylRUaW9eS2AxMd7eymcrE+7tOnfpvttiCddC0jXVdmlHmbQPu
OmnbJUHpwC3I2hU/A6fggmQb6wQP15ogd+FlW2FBjVnG2D/bv2DjhwfyL3XXeVoX
Lm6BZ2eMLFZExoescSW6U2qB/qanglcNk/s+M0I0EfZXe7UoMAGcuEISNv/izEk7
cLTLI2HGHbw5chE8WZ3Uybo7uwzf3RzCnHAc9I2Yf/v1ZHiUFfsQdty3BnqvyA4l
EgAC204plrDngrt0PY+q7LCf4TH9893wS+HcLzEhGc2yKmCzWP9smNbgJsqM+NGQ
bOtvl52qih/XU/42bsaFN0IRRKJHfVcUV2g4ABF84PDlmQvDF8PBCcX3Re07Fofe
5p60bAstiq/0ZxiBUCNKBZ8Xi7+NSdS7GfL1bE5qIMRgeS7MP19Gu0M7ssTGsn+f
gtPxaImmz+jgjIV3aGc6UA3nrcB/h+zMl1cTX+rIIJ3zxcc7Ul+Dz1SIc5TLtfy6
xknU1NAhs+O4eHiJ1SiQk5nRtoQYig6wL4VTGNBM+6Sm2OQSDccvyPPYLBVWpN38
TYXUJ0hyegsqm8YiphSkLmJVeJjpLFef1G9bsh3lCHj+DJXHUJVrfbphdQk4dINQ
pDoYIe3P5L5zeM77x8EpRZ8USXn4hYLgQUU7np9xhizVVYMUdUbDBQkG5wGVgpju
2qIl9+Af7xemEWy42stc66UGWnXAnqThuQYhtV1DCzNwifMptIZekUVlxcxhozhz
Fc0kEAFrpzoPjR5rvTgdmqSUYtJt/fpgCIycVdzvxA9CqPppmGfpbe1Eqy/WBBoT
TlpnM3ZM0Fp/TrhAF0vyjTCxUFBMIL0iLxS2NpdpYk6O6KYWHIAr7MfPohuJDZJ3
A6Ee2HOd1EmrxCr+cTuAswn+KPssL/rSaONrDayZd8QLVALEYmvdM796aEV1fTLR
8cUgUFqWpc0HFW2OA8287MnhDbj432dwmKZHBADf3jgsL7+qLdTwqr8Ht1Da8ktI
VQohUy3D87hZEg0302wLEdi4Shi2L/Yo9Achw577rrxeBe0ffXEuqreF8pkZp6gx
OQMG+JiPU5k+NZtaoYOmTRLtfyChpG7zoNNWyRq/PA6aTAkCjrn0of5NcWRqUwdk
LzCv/ACApvlWq152PzENqraD/8VGJPvZ6iWLseJBHnnafhQQVFilHtWwDlWIuRQi
OMHfTgzhL6WzmhehjCCqPjMAEE3ldswUY3JC6ptHttTF7OuMyLzIJQ/p85P1Os34
qWPRv2EDQ9YhWswlhi86TsCU3nKN7D+LXejp+5AyXt1YLChwo3KRyRiz8AJKDwzC
NGuXuOK51zPHLUlmTBDl73sbWJHOjgMOX2oBobOnaRSL5R0eH3TnOZbYpQ125HSS
DyE2JG+QbjDRJmcRDqshFjaLoJQwogb2c9suuDCB/Q8KwhcaBCHpunlPqeCnFylD
haU8SP5Bztw8c+DAdOu5HENWNVj0/wnYdHzZga1ZjkRwtqjGR0g5saKq0PiUa1Px
RNDeGVAQ1xor+fkJaF92oWPZuqLa/vq067XJBwCScwSUASUPz1cwnqR8If5dHyQ7
kZiXRV4Pyrqq0F9FlXC8DYBI++UYfhsnE68dQ12u47eSg2KAclxaOQ3D8o21c61Y
2mgaS7ByTR7fYYF0iHfGpCRkl2dTfbDeXxyK1q/qTU1bCKg8xS7z/EwQz/1siBx4
tGJAgf2Yf8KnfD8okOQaMxQVWdxlxSosZ5+LjS1XqQC43iLOStbxTDoZJnu0lPuY
w0SAYeOGhudP4IY2zHnkFeAc9oLO9Mg5zFNG0c0jVHjj+CMHrQ/EzKBaDt9xTp3H
uSJog7iAAcMAPHCHQxjyf/XJlQveBQGFxUwFOc0LUDQw5FZh/l9Ob5FZrerxuBvy
DwHmJsjiO9VGYxWOi1D/5LcePbWTfI0HViCOocEnAlNiu9IqKFEFTzVDyVyTMtL7
U/qKRlkWX3K6oakTr1osr9FlKjjpt+3vSXJODRN2L0BMt2a1s4ZG/4zcOGU+VNgs
/mAzBbPvnnQGO8+lJXiZVfd7QGBefNpuEfbVfgHnTKXHcfMJNP6Zj4dkXOsYx2Sx
Uosf/VN9Zn/FQ6igf2Eq6oKsGzEF87I5/7Gu6gViXiv7Wy4Q/8Jt5RVidlKyDR2L
QpjTW4ByX+vtt1vS08vQIccX1CVoZKMHtgsJd+zN2i7n5gtXkB8gJxbXP9VUOJFm
wBUl633dLh0/Dx9hM+oNJjdBq/4O8iFOfSxlCxIxz3xwkQL/wor8vu5XL043a9gf
ZJUx9xUfIATF4SZPigw92te5J2CvDjUQea5BH0icH63bBta1EhK+lh1eZCZ3z9EM
z9EqVqcaxr75TfTfgyy/yRSg1GsUEiQcs01lQChOv8RHPd1swupl54xutzMnKTz9
r5khpyZDoxgJdhDxk05PTivrM0s9QrtGM+peIZi4a7/xHGEHLp6r+7PNZ3q3bccp
F/lxLeYuN4EVwapbwPVV8yHZBg1f5lTFKRVsekaWoG4AucxyiehGh9jGI7CcBlxQ
XY5/za4mvJZa/QeVPpk1KisOTo+3ortoPhda+i1xE1uu78XlYhvXP1YqQO3BVxEl
gH7yY67qHfYUKA8b1awMyHnLrLQXlCYHBk3OkfEGIBFOzQEAJVR0aTem+RVAgdsO
XPEiOuitQCjbxohcSgk/dFiEWY25AvwTUMEc+uI+jaxK3x8gzPiPCaixeZnOFfRi
fpfNOUPmymDd2hpoGpe/mzN3WisuXwQ0ed29mzgyk7ZKcOU07j/E6RBrM0lJTq0Q
ko+GkHFj2lcFUrWd+ZnjOBbuoNAxFmUajuDabi3bNt1Eodn/4TnYXhOFCkkv+RXP
B3vsPF8EiL8+cZA+3pOduoecxFI7c2PWjD5kFcj2Trc6/PHgKteqUuXUpu4OP89Q
N0Fxp7GFF8Z6OX2CrNL6u7LA5b0KKUMJw9vMI0rZPStsB5JbFmQpPO0oJ8vA2QeT
6dHVSz3oVHbqQMwjWa4mbYwJNNywq9jkgxuD8oyPnP1yndqj3kr3iYBz3TOaXFtJ
EccwKzyUxtqIR78Rgat8PlPIeoWFXw0clqr9VdQiuEwDMIhzRygKOEWiGkkhnGdB
WH9h0mdx/8ZPWUnORfvBg6uID53YFGidMugt5VTDs7VZPpmFRPOsRLZu8hS3MRhA
brTVB5W2dkOeVry8cL1vQRJbzlHZuAKjdD06F7mVkMXnIf8/GXZDxjyTCU+Vg8uR
mc5etmWjn//nwFcVx8ixE9jR359ExF7kydFoRvmo7qP1zh909G1n5eBXuEaFSXOA
F8zL2FH95z22QVRCND0pVYdy2j76Ws5xgwClz2/ponkYoc7BXm4bZJlVeYzKPcxB
m5khSps/CLpCUjkqYo4Bs2Z+TRRDZpVXEr5OYyOn6gnBpnuduc/nQhnJXsCnMoiS
4dCYi2LvgfdCol/uoI/a2JwJtdqTH2h35WUyIKlgnvczLBawzlaBPZBsqZwerqBi
o+EghNZs/qfUP4ijHQ6I184CpPDUMfl2i6fPP5egYR4U9jJQLQfIF3YM1PFQS7iO
kHK7DApBU38xeYFRgPNsViRioPGelQ8loLmsoUlKZfM6s74xRS2M2VzX0cc7uK4Y
1RETAT7sk2hp2uGMUG+yo8yAQYNv/A1EERnZCuNDw5NEMPR++vQWIli9WIw4VeU/
s5ERUDaV9xZ1WtDaQfjZg/MuRojYuNH3JaW+C46qkijG3JLsUkJ310KNkXB1vh7R
bmG74a/jvmXTnGzfcAEbOG4YBGAemYXSB7Me2KTZjogGBjUi0xp/5ciXCwe9oxnS
yDLJjtf3gFxU3QvxKKp/L44mS1bedEH5lbe+vO7ahg0yaCIV4TPLrMe9MCZIpwcg
UUnaqmpTS4058mRW+lyH7hUxV2aoIUp/mgqqlYFVNkhmovbNvkTouxYGQmq2Q3qD
+Uc2sQuonWGV4RD50PnHqG3Sld20pBt0rMWPw6sdGFa1mI0+5/gVppaG1b9LOEr8
fdZ/JwolpMPgGTFFDg2Bf1mHIgHKPwZe2wYAfbvrA4MPqvKKp53bobmXqxBf0rvJ
aUE0yWEDhho7H/WeS98KmHAZopN0i7aumHLls5Y/SH51C+G8IBRM1KwWxD17DUSu
MAmww1N7DH2TL+0XyUyV8SXfm3gcVzqblsMEACBHh6KpD7S8tvPfSlwVpXQMlYMG
5DATdECodinB0iCO2V6htFfuwKqsUDL3JRQNa8Z4q3sM1baFuasiSl6wFelfsQna
8tXyIiiFhCRbWnBZr8gUF+GSkHZOuk4fFizEZt3QKy1SDxXMATHKvQnAJEVUQRyt
GPIkiEicFIUSQP0lrC7mSJPzUcnwtfMTgqHqVNZerCyV/qP74wpT/arl9cI+LCl5
Lw4yM70Mfwm112eZyGo1HgMtnGsE+ghfrt0RCEfauSbVx80bfzrqadCZ/4GfGXt1
kJjN00MKfqS6TnaE6WAfhhgzgWK/NKVpJ3NRnRXhhasIGem/WsGUC0+DGtbmdEUj
no+uJOkDLGfcyLk+xzhTU+UC5fDuJop0yaULppIQqCzTvDx2Pov6KHc22W+fnM3Y
kNtOwd4dn2bdYXDQAbO08NAOv5q+u7+q8k/Am3ZWzG4R/C3JyWb8/PO+D941gwU2
1N/rl6O8v/bF/5nk4fZEzLHeQmy7e1j3k/uIlMOY7PRLXj4ZbKN1akj5jeYxCwQL
EY46PwwNLWeLEBSuNABT4VqFqgMzJtp/DN6aec8MdrVK8OJYa3GbAoIgNJo6RQ12
9Qv3toGsv3KclQW2VcgKonItZKi4Pa7qMZLObfLPNEWzP3RpEgq+m0MfwtfFTnHm
Gq8Nx6tKOqjAjDegOlCf5FjkHaCka4fnqtvKIFSm9Q52PlA1Xa/2hFQdfTR1iqGk
o5ygpD4JgOnK8HDgn2knmh2gsG/CiEP/mnwvjOFET+IWeuIxuJF4jpd/isQSB2fu
WolZej5lIFNZej4IKeFovaD06i8MEiObIIU1/cuAeZa2lBrqkf8Krhzk9RNe470s
RROc8nK/UI8mLCK59Qi6ouLdYR3SmyqM1WBPUo4wXBn2rti2YVZuamTYK7tMToZ6
4+jVGn7Os5Zq/BX6FO7oWw38WPQFm33ulB9uYTlBFxwveUjIhtg3dYHM1BYLxEg3
9T6T31mwe1bHHq+fwiikwhpThbFABLQcQvb5Xc/JhRnGAgS81aq3+OeYauywKFXJ
kRIAypi6U6msTETjX3YXS1oqOD9Qv0ThnQy6eohc7PU9GWXwsVNplZpq8qLezV2v
AFdT3zVs232Vnm4oCtA86E7vAJV8sV+8LPXX2r1puE1DmxC9WZ1qE7LugrXXX1gc
9zmOP0pOfxdBpeZfa8m172bDPr9LX4IoszXM5YHnuEfYNnaCCshgnKtghQypW9uS
38gURbZVpteG5rXjijhEcy+txmKDCH0h19e3ZqO2DB+pl4LtZu8lrEeDmUtNzgwd
E5cTUQkPbq/9YZsWNw9Xy/ySBc0Wj+InJhEWEMLP13X49L5AKdevA4NLZKeijR15
xNBq9xyJzAJPlr/KvFdIc+iTOGXkf7+fR9DI58yCBC8YmR4Wn1oKQKDjqd8JzgLS
2MFgd4nVptrAq6klhjl2zlOpZ4MTrCu/9Oug21+570zCv6g57raH6lp4DJb++0Kj
gjm6F504GmHU3MUBtnvaCvp37revuJ8/Vxpt+JnAMLqsH6MeOd1c3hoFLhgORYHT
9asIyLwKDoK2oxp6nHqIbkpJ+9WoiJa/DOGlMhLJnHKYLaSaEhfQNkgJlmwaZqYR
ytBVaDSwXf05jzrzsQaBkEA/2JgpmzlxdzDmDM4QwGJ+ZMSfX1XtVhd2nsUyzmVs
HlO2p77LL8woKERKPY30XzcNFxHQLMDSKxi1ZfEshM9w11AQ10xmndyw7S/5Y/Bl
QxcjkdkyqNfmsYpEv6ZI9FHxWFf9BAc2K3r6OtwmCwQoanJBWQCqQrEz2Hezah3e
346CbOYnGitvkJhYIl09JUCdb8r8/fszyxXlvnnRBkpnWPnbAJ3deY6H0uIDla8d
N1Ixri/yn7Caga+L8k384B+tpG6qDEquTA7mTRRAxI1qK0pnUjInUjO7bXVjw281
XNu8slz6T2my8bUctnAMUYK4fYGJxl9xh5ayiPV5FC9cLaqwwSH1cAkary4FeRWf
QR8weltn6jkOrx74iSRMsoipSinc3aCElbqu4t4IRKNs4EInTIwUWZO7WtUWN3bL
TikXbbMzLDZIsB+kAl+f6CP2cTAbi06iN2A2awkj8pSm1Q4NUsA+gPw+vUowiWi+
k/U8OCq9kh0pWBpFdDLlXMwDqBf6jcgw9ICz6VBMy5Djre0HsCmVooNbCQpgkW+5
Iw2SWqnX2QMEET9wnO05BPA1EZewb51h/vmahzgmyB+9n+QAgvuUqIAaoKeCK5B7
MQcMapTu5j4+xipD4zC23MdfkWe7OR8AAiw4jHS/nnxgYQY8fmzoUertN1OOCW4q
n7WZM/JXQv0WXx8wNNMDJNAINbjtQmrRucs7CAWR0QjFS3BgQIhP+mOmEtUFY8L6
UgKGsULyL0CGSiz2x3s3oIGdmbPDKzScBaXXipcLfgC+G6uuH4QSpSTCYbJ1qtb2
WbcJ9V7FMSXts1XuSTLoaHwrm0PjLY/l1Cvi+a1BauRkU1WX/91ykV0E71iDN17J
tAg/jKH7RSxfasZPIM6M82ZfS6a4DoXcgFgjf6LSZhrRkoFxb/sgJ9dV0WbbvKEs
3rDQLDQqlZZ7eSzSJbICyrv93qAX1FPQTRQYaXkw+zQNj20FRhYMtsYYwu5MtZAI
qp8yEV1+zEXCysYZh5pGUPUTrsE31fwDrdhUId62AbAxZH4ouiQUPgyrpSJHS4MY
tPneg6etEvhfgL1nLO6SHt+utH6QkUyXtHgWMBkfuWzTUtk/akT7SQCDWOcMH5H4
bVq1jl6omR1YF4FDFpLArB/J5jDmsmMsnLnVln1hw8qBCjPk6oeXN2YzrlVbARyM
nab+N53ijHPFPUbq0cgFdm5L324+l+VENpk5Nr8Zuw4mA10UFARZUx7/OxQ3XvQL
9NqhFo/0CtjObrAJx2/WmZygKpb8lOuRT2BRRZSnPKUfDRmOcEo7EHm7XfesJnBO
f1YDT6KksDTs1ksa5Qjc+jyZ3X7aQ0YB/wmwY7+AMur9EYEW04ix7cZ87x6GVWIf
XrRjHR5wCkrT2ik5PprdX6R58CnRhohXyxBXE5CgOOyXRG1vGbkjyNhxcuNm1hCM
zbpoTI1Dwb/7HjGDSM5Qhj2pKm3i5VSeWvOQjzkAnZE5KznD86FYNs3fz9gH/fwM
EgK/u0T3iam2gR96FiJu1L8DT9eujeptY/T7J8wuqcrwKYTij1FGmYqGM53BngPB
wNK/pJQLqUlQXn9dgt5rFLAVINMLpU/zinYHetHubA73O1O8Mo74XjbegCtb9XZs
Yq+jWG57JRNPZHk8vUmmHdKR5lyxfwSaNSAmVWtG2RL1D9biBjivD3diy+g9FFNh
efFFUyMG70SX8p3YgDvTBhPgzP3rRNUICnCGHmKjadMjP5R2GZ4mLT0VPsF8gHCE
ag6Utk+N/Ab0ERL6NO+yD61wZMeGxD5nWkhDQfDsgszLckZExZKAngzhXgpItwGn
g36Eo48cBSqkRPl6CgiW1l8r7+BGnRR/tEhyQ5xNrmu06G+fN93s2tk4ainru23m
SfGGEr9S5CjoZYSLko7Jq8vLNYCOo69PuF33QgseiFlUDevQJTdcTBldvF+yXZRF
xt6ivq/ykM6GZUWdPaKf0yfx+KyYavYMox/fR7byrljOLi7tVOp5KHYGBH5KdzTj
OD794WpJsRTECxGFbOO8APDJqp7sHJIG35MU7Yf8sKipiavWuyw7bMSZAP0BkgLK
KN0oqnBm8B5FplMs9A9EvaeCl0dEJJYLPZe9htm8J0aGOkqxZsi3jGp58BKcCar2
qCyspf+pad6cWYqSpIzp+mI93HbzrkBdoUKMaxG+geG+/DhLhVFgyW5i/C4WhST8
f4vBbYx4TZ8uv0o4CSmvkdNQJeF8bK2o/ATz+5YJBl9i51v0gxZu5ic8WVcVatzV
zV1NaDq7hAnGbY9byNU8RiODCo/CqX6fUtfy2r21N9f0O6UZStCowZXwgQ1yKDt3
bQe/YFXcm38tXA41+6RNydu8u+dK5Hi9Bxd66gPZIiq2RS2/smSqC3bcNB2/AfDx
vadlfM8uXP/KXZEd4CNkugS8N3uvcLyw5fZKK05pzbfGGEPweSSG9Jxtp8c0qgQo
DznMXvvVbWsFDzGAX42/ug5p+l8JJOWM+aRY6QlWDLWYcoVt5xgeiq2tj79/XQi2
in5MskZlW3jOxfGv8/9Ube5umKs6fUbq9v8R3xQFFN3rMg5LU3CY03vErG/zhHCs
iTeCLUPlrkYdQ4hjHBnW7pk+zd6RwCA45B/Zx/pF2U+pFbiOmYmEdqryiolyibW3
YTiQRR4dUxqxCAzwR1SkIkgR0W/deDZxikGf36V1xamLGTHG4TAvBvCoyxC5FXXh
idxxVeseO429D/7Tm6UvmrAfjpcuK0pyNu7Wzlb/Z79GLnw8yfPEZIjoW5ISnYbR
muiLDefuQI8GfhHZa4mkAgusKaMgR20bIFaJAdkGexVy8CryrkhTLOEoksvrmZFc
zklIx8uZWs9mQuO0gh3cN87xrK44e1bcVQdy1KinUPPAlDBUCNFo7wQ1befOVb0R
jYvYbW5XXlGlBMHcS8PCOIEmT2+DeMQ72tO7zFDIa9wm26z4qmnW1fz7gKXIWEze
9IJEqbjleSBmivLLMeWPGA7poMxOFdPiz10RHU92Yz8KDFoHqQDgK00Ak3yA6KLg
CgHTRf+fFI8mISww3+YGfOd7hnOr91cAK9WXNFmR8nu+yc7RK//XJWfbUS/7pppy
WeisxMUDR7JxVNnfsJi7fHURETMyBM8uugABXJTm8ZP1+SOn6OSudQbKejgYMHk3
k8TPJ4Y3NVgq4mRrWIN7edd3QZluy7VL0zL66Lx+aig3TPyQcTnr6FklPBDjykCz
Ww+BPLeqM86VKa/c7J8H6olVw+HcD2sLG5yip6mOnzTjucQ6b3AFdNeVQr+E0dD7
LJMgVQkI37M37beg2YGbl/3CvxpJiqnmlATgpCC1QPr0zmlbi95XrVCi26IZDoJ5
kiiFa50nBweBkVo2SLIRLyRYnXHNTMyoqhaujm7vFrPCgc0HwkyV5eXNQ/GHiMoF
aju3P+UFv10VQBH3PcDY4coKEpX+4RqpIRM9afSYmtfPIPz4UAgC4FN23lqIBjI3
QXm7G8cPIZ2Ih4muYrEOfXBKMHz8vMtGkHJWS72kgWtwnkWEpxkZzrpR2Jeh3dn9
nuX4t/2ZLE5tIDKrJ5M5JI0euGHBU3cto7sZnLCu9ausBh6H9jUn3v1G9F+5Iw1X
rDkAKKShPbenDmnWF+GYWN14g6d0KQT1gdf5qStPofAA6KTinj78siP5/VV8EZx2
mPd8XNKyLTbH2QqudvtGu9tOm1YGM+BbvtQU7QSU2hWoZUTzw9LvLxhUJ/6VfIGc
+6QWE+r/t6m38N2N8XPDMganzJLn5d3pltNZA8KAqiL/M1mqei0RhIywr7c/B1Oy
YIZpvBeeceJBsHneez4Xx7BDWh9l7zTMuEd7JmQ2pD3W5P5H/lPb2WVyer4lOJrW
1Y+H/sDOq9HMtzQZpLGgrAFobMLSlq4CsF1OoHxS8kAdBsXdtz4X2eZkNMxWNUBK
/6QxHLrhAftA8neXd9dHLRj3XtElMxGRMnPvn0ZtxyDxmMxvUHXZg6K6snrCXYD7
rgI7x92yGayEI8+pLhCGbHMQeZD2qX8ztzjiDGUAdyTPGZqunzYe0QYEq2QTZcR/
5jI+j2UR8f8sftYK9h3bIiYCBDGh8H1dRD3eM8rVk/gstuFrmDMddNND6HUmM9rI
ZYz0Ty3hUqQVvgCTR7ppoWquXuHp9fCGvTciQOb6jqQK2ZFLZ2ujYJgHm9OYueH/
wn17T58rjYk9PQYCBoIuFtxjEluIzd6E7wz1DJgVRPmm/VPCpLT/pbbRj5fUoG+p
sHJO2yYoDz/qISCRbpbI7EJ/W7wYQ3Lc+qBn7TAf/O6ukjjOnSQ7elXxls7e1q+c
oKpNjAESniDxdIlqulUWeIIht5U8qRbQJxSsWjJVVD8E7YEnuF+De+llTgwP34Xv
s8QccDSR15Y+uRcUmQhQjkE/WIP/PlhdagXQn56kKTg4MRY0o8ZGn2rOEBcKlUJ+
RXPdPAJXn0RQmGUl1kqPcPGkF/WPGGQCjf+mlMpPR5fZATf42XiRTJANUG9tQYNJ
ZlGXzgyd2q8W7tdvB2aOmmyBazw8WFKjZdkbyGwiLN774/B7vP0qaE6xD2nbNrv9
M6QHu35Mjp8apGkGHgJm4T1DATlxB2LmXr2uvmULiIPwTgO1leV96XeIlHQ6UIYj
D/JTq6rZWNFDmGROhkbFjBl3R3LoGSlwTcgcNbhp4aEZq7eDzAPG81iwg+xhghVP
bayX1cr0qsGdepajdNch9VYDzJ8H6bMr16ipHTc/w4oSMQtBxZxbmrEjsiexhbZi
3/k6j75oPjh3+P8Hzaq0oMxAO6zsDXVDu1zKx8GWMvdCap8weecUUf3R8a7sdi4e
8RUVhHug41A9YZZBYdYNYTmzx+K7jdkF4Qt7PGyFMK0oGq9rSLCS2QGpQXOyEngW
PgcnNSFEfGHUaEeBF8qu0f029zxnIOXFvViRDjLL96O1vxOgnl6UnFBT/BZk2VjQ
P82+KvLSqPDOhe8ICpF4aSeQmGt7vS1C3pdFJJZgWTGLX4Jhnd4Y7gIBTQlmGY/2
KpGoAXCBYmatnHdnWYIPHKYBqlQpMrr6NR8lhQ7CLW7qB5tmmDGgITvg+5zOt5p/
GUUZmZMl8sDSB29Fv7CRno2Z+r428tmLo+A8IVbdPxDvJsY4EgvTAgcbGVu3IfwI
a59ktHeBnrjijghNfwn6Ztv/8DYIfDBzVsxNpxZSNRdDGt7h9yV+g566o04K+QxV
mBC2xJ8gtiWRu1eit4jjPqfoCgwNE676Vfyk5HvVSgvch+U0Ucj5xQv/j8ku8Dap
IWeX+vn1Hjg6omgZ9sbl7JORPaxeqzZSjowQ19QoKLP2u6YhwLUjt5Jc9sK60PDi
0281YYqrO+rS67CYt8ggT32lDMDkKz7bWdOOnDwRBP6pacDQNBq3E8Tc6MA58U4C
jw7diwe9dXIexRlXfbIoL04ICu7nrdP66crsNFG3iZDcmeGfOCcsCXi2t0gi9Xbj
nVwc2e0jzHI3pmBQ44eCjSX1X56NAIUo5XTfuoya1z5JUCQJfdqnLFMjHa2t0k0r
RI7Uf9ngMkPlKIujZN71jDRnc6Aiuj7A4SxU4dI+0/8tSY3Jy9Ov/1pvMwfIXN7e
+GtqToHXkAn7nbF8sxXaSejQ6Il+r3iVroT9mBCODBZtpdGSPxZa9U6S5PRw/NQt
zUD58v8Odhef5SmAG0hIyzMTl3hFd+GvF3OoPKqMRQGeK8ukIqOf4abGjwZdLJZA
v8x8Q5MhN6T9L7psQ7oXoPSlwj4Y8Fub8kCtrdfdUoIUATlQT7RbuYHlyjnisrv2
7u8gx3tvKtPOa3jIp2wNIPrcUTNBX7kyJMyZf8SfSYoWjQjLwZAjD1/eEBpiYIos
jAl29g1iwLsQAGt6HFa2eHjlsvLdmQ+vCRBdyn3AgIt3qOBSjVNTujf+4Vf0ZRFb
9AQf5ro4bxOUD4Tr4LW0fn6MmXAzM3HPrZUuDciQ0YaNSnEV9kCSYip0JOWbF+UD
QvG03K4j0vzbfjJTeLJl00n67i24Pqz0K5QA8oo6cLiyLECTKrBwtRtcCfmRfOhm
vs7vAsiyaA9HhG+jl9khA1VL2Gwt9aOK8j8uHOtUwbC5tz5pR4dhevOJmITI2m2h
DEci9NpC8p7vJWYymQXeyTs6Z0a3AmHyUFOgToWvWmYrQ5WIeFW59+QvMXs1sYJ9
HivnLEG8VQHtM0p6SjiTso9iYoSxGDg81WjgnBlNhf/Ab5LWdZaBikLV0rKUpelf
6WoW9S7SYyteootCjSpN8bmG+/brnZ0PhUOAfWPttfwCl89Ri3+9+QhWUZQy4WXx
U7xJU+wm+QUpbKZWaWJ/NaTEdDBPinJRMCo2i4bYV4sV7ifOLxMizVH7LDmBODMl
N12UYh5w8cZ+Tvc85AQ00cbiessvQdzWmjxwFk8BIZ6orUii1+Y81oNIeCCihKqU
7BzbbgZCkIsaYNvbOFQAAtp/ndy0M8/JSisHzH9C4aKjGod1e6wGYJRPXmc+r5AA
/xMVuhCue9etYT6rYsPHstOe0YAEl35fMZpbiVSrAVCxVM5zNKbfkxFUBk4gaW4E
X5arTIsELFrb0es1s5WMrxpQFEkTEn9ykJraOiGtwJ6g44ily+skhv3lO9aV2/N+
zyipP1JlOmYygJODaroxbRu6QMVNyq2A+cneHeZKDookicHCNpgDqqp1AdHkmmww
9E0tQdSpL8ZAUd5uICyje6/+LGOxxUYE1UMh2obx9Wi4G00sGrk+4SmDDmPpWzbg
1JvPSU+xjyec6qsRlFO1bm5P32KGWa6ObUO1mQiw/ysZCHZsR2L63LiLJPrTBTH1
wkq3R1WmD+QAUaKnKF4dcGQ9ToYKLNgzppBi2qdTRhp1y2at44ylK+mn7YR/Dme9
+c3LIfCDp2f3z7+ie7y0kM8Sysh/YG/Wf7we3kLrZfdGXiZ8BPONmR61V4vZvJpZ
nTerTBD7eN//y7ujimPMNAFD01YCrLLxeFuOnnByj6/dDdPvtdx/ibW6gtHIbojd
an2u3yL2RRhdQ5VQn1+Q2kQ6BhwsuwYCC3oVIKd3M+CNRnQvI2HDFdlyQ/5ozk6s
RpTGzCGowucwzc7lcxuATszbmjhwEysCdHyccpgz3VxDldWwIo3CwWDZzoh4bODM
Bywg5d++BvgOhdV+GuLj2RsrtIYNqtBvpR0K8qdVMjRGf5IsvkwT2WLyfgZ0gGec
fA0aQXe41XVLvBeGRD0T+VMq1N7/Cyv95rtyu7vnQuou1FTEpfRGdDZPlk3VzVlI
G65HhN071O+KOG0at/oCX8RjKB9D9ekZyTnnxN6KEzDTSja5QMVRThkumCLLHn0X
Dz7yhFMtJqcKTIp9u5XTXsFHeX/ZWAzB8oX7e0CLyx4xHjn2E2aVUbXn0DWPJ+7S
zbT/IpudQ54mkfLnGxcmk1oE6IhqyhJJo+zZ024bai2K6Ybp04+bYKTC0D9RbiiO
1cLkArmWRpdITlv/ueJwiPH4PAFTKMFZ2/BWRoGnZ4IUQGaMRFqYMzhQaQ5JCY1d
tF6i2BjMaIRpHwUUhScIJdzbZTFXZ3yX0CwiqR79r1leI11v67aj3JhWnzd5Orwb
vs706Sv2Iy5FLK2frtqzQkU5xWYziqyicr+nDqq77U46z4EZEbutJD2mWr1mkPhp
bF/8rLjhSTs/LEM9guJtZaWSOJPOLXz7sDY7m5EEhmvZxmEHJWZXY1cwaALqT1eG
CaD75jXv75IerRLlyA730dhkNum53KgAlHBx9QSD34ENDrwtgJSwBp8ckX/vpmZc
NnMdSAg7wZBCH1dPBEwxlWMzgOnTdP3OtPFaJ0f0JO8OU92i3oGs1BqFqL9Av9/t
WdhOwQw6XWSi7Ruzpqx7wHKGTOcWk+tYsM+y9wmBjnVUgHveIo7jjcM6butWRuB8
AvgvvOVCpO2hloUyF5gh9guYXO1tLHpCIbyPaLPaOo8Pge2GYrbGB+e64yfdD0fg
RUOlDQWEmVwkqFDMgAxx4LGgnhKSrFQrzmq5wxf/301lFOX9wcZ2syC+plLSmQbd
MYSK2ICUkK7lvpnmfVwPuswP3+V1yakC9xf0DFFHzUAo/UfSYiSrtNU+6xvaEG2N
BBMV6J0yRTxamVB1QU4dKRaP1oFRh7Ov7TsPIUeV9DnkaXygvHfwGViYgbxL7AMP
ori0qVoT5Q+Prg7KvWWDzHOy0jGeV23TTMpi/gVzs4VCzkKLcFA59/aDgR8DAZPm
5onq+KK6QKrH4spMZHvC6wz8t5QYf09QCuGT9ta7sLTrv6KrfX3+T6UyTTV/kafK
ijFDX3O0LG05BF8naVOoqbJtjNbMfK4tDM1+slVJIo6uCW17hQt1pWUq/lbJy6oR
KbR766LThGYbVpoA7J+AnZ+BOPWlni+ne4cMg9pJdWuVWRwshcUq2HNevKDczSwE
2PjeKirH4TbpoSoN7FOFmX2SDyaFpoMrw+Lt1Nc/yV0P2gNKQGZoKCMAK6OT5NkR
ai0SHGXw6+N6VtTMFUQlzA0ZaJkRttU/7iKdakHGt4+cM7ReuvU2Sa7gNWBv08Zr
6CY3Gwfbj3nyIpWNdPI5cI3A1SI2JzItTkOQHmCx4XM4F0tKcy/wsVuK0rjpqu3+
WtnQq1M+ZOjE14DM29cva8aISl/rK9alKvmgAr8xWn5tS7O4h41NpXPmInbzBMF8
zMRLSh6uS2EwgaTMlFwqOpzl5zNrQ2yl/yCdcUQW5inCWr7N37iUql/h5uXnD7g2
nWeTDllM+tmRw4rvVPcm8OaEKo23SqOkhDTUQE7SqBpSheJ/feODa1Pe2s4CSqOr
eOTg355z1JIibjulUE3FDzIWYIfHQvgywWCBKg1jgr9nvRS96UHcbf91lS4r4OLr
qqeOkEWjyzTgmSR4cgvJj5hU37Ld8cI6CBsmAqLoSqn1oMGidT3/7BeH4kyCQfM/
J+Y9T8YUXJjLoiieb6qpL1S4tZ/rcmGUsQFKNYQeJkdf6VVAC/oMKWBDh2PkHhge
Cx6Uitl/Nh3ulMi1NIJMvxlPrzHNB4t8jh++n7WxMCBnnw0phxG6eAj11AsCJL9b
T34q5afaX1khXuliV3oK0IXzMg4xNKIx56SYuTQZvIPHaxn3HZDS/tiSlA+CFH/5
NkaUkDM90tFLAJId3L3hcVlNwrk2pgnLuwYHS583/35XnWLLi1Cz7QP0l4rdXsNP
o8OKR26hV0tGRmEMrF7YcKriEQ604upY1bmd/Jfg4tlD4qZoAUalEIBYsoProG1x
VyWm+rmCwrdF2S4CeesFrpTElAYp2O/kCha6SMlM08A1+A9pa4wHVgYVb5+zY/tp
XFI0dMfArJOd5Q5SoMMTbKjeAIfZx3Ln/V8X8+ydvjWEaRhDsd03RQnCiSOL4e3N
MDBf4OqoERc3wPSkQdX2Jy3ncFVdRYgIPa+bF1AtzOvyBue10Sj1oRNQBDU2+KB7
ovmMAXXwvfCd6uY5ytle+S/p0FOAgUqOpKZBHH9bY3jArox4HlvPBLf8kFDRsT4v
KxHluh20KV4Nwy5X81AkOM/TjQ0KHKW2DtOqNVBJHY6zXUvbP76xw7IxRF3AaJVS
sfh8/elMkO1UjEQvG/sHk7Dwm239K4JP7N7k5aE7YapT3JCcbT7QzzuAX0Djm1AD
gjtOAo9qwHBJoAJBG6zBjKE1dCqgFPIhdUS9FkvVBz284wQEDdsqaGslI66Fq+9x
RjdFCKI6RoXoTTZrRrKzYuubc6oK56ejF6J7VdSOb07RLhqUb8lRXnFx6dHFnFU8
nLYmIpyPbEZLpBZAYEDRHXcFU1tBQKIWGQPvHsyy9eEOjMWkAOamV6HYn24NV+GA
xpisdPtEVD766dZ/TbrW4DbgrSwOaT1M20OHsV2MuHU9PFhQczAnR9xjpby9fOb5
QhcLy52N3TKITsLQBXAL/Lfm5x9jD0HS0gABLXh6q1qzI32eviuXZV3erM7KomOx
lmWzN1v/QfAsjgLwOARqWV0B1E6yKboDujc2x/MWBeupAE/CUymJorhfZp0cGWLc
HsZxrMpOsJKurf1AT5bgtvwi3l8XXG60zhs8zUyJMzmat5Sc6DkZKndX8tQ7T6i8
QxldzgHoybgra2zgAMVOF6EQW/MmhrzdsWyzEAeWVqRHKUl1HFCMfVN/+H24Lgee
tChLYcLsDHaVMr64z4CTar64s8o0/thqR8F9P1QQxqBR2DxdfZcIUKu6qZQ72+pd
ANe9U23cFJ+AzttUtbIxNegpj/pGkYTS6HdBV4CONG+KE8cFedGRp9AK5b/7NE7K
OAceJ/yRm9LDx8xG4BwsVuds1tLx3k90anPj3YCT9tSxl3pzGooKWgzpNtAj+ZwP
w/+FJV1KOAgc3sVeFKfnz1NlCew3LOejWkJv5Fd0oX0WXml0rU/8iHpvAHBAIbuC
xvkhcZu+rQpMPD8onr8TMUjqL8dkA+V2lyNTQ+/7gsivDaVlqwwTqA7w36MJ4dQP
MwYnx8eAI7XLJqJJqe3+ohOHhObEHsdxxCjR3FS+5k49UIOYGCTAu5UCQiYFtvhX
/AYYqY8kewf1FthQOIoSfUcUu+TuEbK1NVaApgBTS222ZwaoGGkvKP4eoR/kfWau
Fj9WOjkEA/JgVjJKR9gvOeF7WG9FXio+4PECavxqny661QfUe+4f6QGymJe8AlsO
QLfso79mtnQQQ++s9yeLJzKDe6zLVxmctIQqJlTz4XZzRcpN1dWdV2PPUo71d3cr
UHzQ0bs2suqvkLVuQn3xN5MtjasizdH4ee816R5kJgZLaeN2ZcK8sBNfPG1hOYOk
1ZUAUBJjVMXxFVio96E0BOLTQ+Cjr2Ccu8XqJHyKx4JU7OhWrxqWDH0xnNxXnNKU
pC3uGCGf4sPYsLjW8IZzOnH7Y1MDGe8TrqZ8gl3L5rkz3FA+YZKMfD9/CBuuFgEv
6ZQCbpCF219jHicXIJuMYaX9KTuJ6kRLKk/1dMLN75BubRDWHEpq9kwdRnvIovrm
kYF3ee85VBAtjsLUVpi6v3WWaEKtPueTNR0J8K2Hq2pwm/RQnMHWj+n9p0MfnhWh
J3k+2PbULknPDmmYKS5HY7BtufdGcv5DejusH9Cm1p6AD/ES599ARqUN7UqxhPyP
5Rx+dqstjSiMxdotIf5BsMFlDYTNA36iQeSHggIF9mtXeb3aDoD8hsd+j2y7FRbU
u8AmJ/U4fbQXfOSuStsoiPKHiOcAGt/sdRcchLrhbgDxHb5QyUP8HkZnYolWbEw7
jmtNNynwgJtGberrHS9ZbYFiCx2rZuuymRrGihaBC615pPIfICN20xAPY2EzOW4N
udUu8yZXmx3hGnVYsdqbVQJVhEzw11NU2Grp0DohpVYfUhfjuGS335ZsNHKXx1uH
1bZ0Hg5fD5XK2z881PG/oSDJqTiyT1caoSXDebIj8dQpY5nhTHyKRIj14WmuFgYd
SfxJCzV09mdV2S2jAJGna5znP6jDXNzRS6BQ1MdBqVMGeRLdxOGO02yA5Yc55UyR
ZWmAbltXc6N9ZqLKpxESrhXzPHUq7loSBq4QGGg6wbaLRQBNb1HEKpKlDtLYOwuu
P6ajEJadMNP0ijclF3TWrTh22vNJHfGtVmqRugdPziCjPhRa7HQJ4o51HXLH4ksZ
eP5QMSdwLpLBHQAoXuPCR36zwUrgxuCieyH2WiZFgGC+r+LUzGF1h+XlAMR0On4f
khO8xuuylxVJl4eXI7jSI1s/Xflz7LsEYyFwTSsRDB10dOreRySKSWecUhBh9qbm
jDD0p+tGhEgOCb68z61PU09/poyZGrjW1KT3PKsRkPLFB+IvmcJ3pssHRe4bJFg4
a65g9mgbJHmBrjT3Rp+qjgflSbATsEFH/xKb85nDrxI8E2z8WHeZsPRp/SB9QHef
6MvM1wM0jxiRIn8d3tyOxexmE2zr9W3Y0xjP36ZVxrPNySZyM5gLFcnE/QBPdVHM
94LlQiDOfQvqTIkozdryakP69cHCPkVO0RWlPinH3ZdXGzbob5+rxLYIRXYmYFf2
oTFmavXCChIHAi3wrgs4Gvh5feMD76qDSegAWKLay3BwrO7a89Rj7T7fiB5j9NjE
FCdjo+a7KNxBvjzVJqIVuXCHbHqgWWOsQOisWcH5EW1JHxMGV33WY4w7DDhBOK9H
P7DA2ewIaA+k5sr/rRlBpnPXdkOuK4S2qnOyQEgHmNhCATEGe/Fn0mjxoJzumAiS
NrShBtxCAGZn8+1brfW1tx196ZEpPiUpXl6U8nyvkxN9oeDN1BoF4/T6HvzMmR0B
12kTZ6uOtN6Xh9/iiWILP85IjoPc206cr0yWnVdwMKD5JRHMLrOHVbfPwzh7ojr/
d0W7ej1WJEz9PYLT8qirkR8rU+BIdO4LmH1FIQyATDlnkGUCz2jUUbWucUdTY1B3
PpC9y8ysQ8wCxFZeuT8HHAwXwzZCMxFzEOXWiMjJX4RXwD71e+6SOWj8TLrMuVGL
yGG+Mp3Xa6KBQuBmSBKabD5gxXyntW1kGcEVFX+mrcECn1zRZRoU6W2T0ML6u4rr
r4oTMVn/kA+bVTx3CTadCCmQg5ZMS1LZHcc0INhvhJfGLqRIUsEuPZEimirFfG20
JbK/XZhnfNkxGT/5/HPQVt/6JZVqQleJIPsC6vPuohJHIGY/E+1gcMfrTB0kV8F3
pgcRfsL8v1njryzst40l7eJIOrptdmqo+M7Zp3IRMIAbZJb93uQzCsqNLTv6/z9y
qhfR2qSE5AIphKZ7veW/479hLSLZy81ZjaTSXJrepdVYMfEukXMjNfsvOGDz1DAi
1O+pSVPm7Kw5fKCNka8fTNWoSooPJTLjl8PkmwvJztWk9gzPJVwPW2TARcYfgN35
6JHcJFj1lvmncbJ7WFoWKCkaRoqJ0UvXpQU0BMIip5rVqq9y0nMCE/oDtxWFmQBV
yLBYrfLlIDTVkwJKfgXAz/cWKlL0/MSHbHwkstKoMs7+X3f3+L/eA49tI+FFfarI
jMIwlAIwLDtnxiPl4ZkGVp44kIvHWvRyW3WoRzgyGPb/4qP//FE649f8UwefdnCY
ae+sPt+yUUChNTBxYXriiLfDI3QOk3jpvpm5mdIqAMuEsYf2voiei8N5YrTJtrZa
EhOqOgueHb0Kc3eF3i3JkZ4BPyx9dP7SLlEGy2jpUQ/RPgtJdFcF0YhmrrTEv567
trQchYO35y5jGb6ziJCy3KsH/8sBGC3fweRZbbLF8cSfNWE54Z6UIn3tDKFDJShO
LaVQHvVr/NKHZo+hyNVNyiecNLc3SEgvFNxdj5j43DNaISUWvMY/OA6FkAzFQxNB
3u14ba2pC3YGEfEk6vtGKleoE4mzdgfp3KqCU+sds9Q2md+cxoy6Yt0ie0JqH9Wk
WQxdMZ2NVpxwe4MrhHbirF2XIIS2KJSQpMarCyWaZDjyYUW/gbpVvINcqx1Hml0g
VA0rh2JcbcZOqAGhr7g0V8KrnrWAy2+09S/3Tokdojv7XkbJkfIxCa5wxmMFTn/Y
vbhmvNmtI4Pz+zIC1wSASpksSdH93fOQDKZSW/yOLF/PE6dcsj5TFBk+nCZ7R9mJ
wV8LcRwE/tAchzuf+44ao3jyTw+IPQBB/+vD8PK6CRnwXL4ICsDaS+z4/pG0e1eN
A123sSt/hrRaIPkH2+cibs3FKb+3sv7Bzv40fLcioUKXa/HRpl6XnbHPmuylX0Nw
Leut4Qm2iaICU/t/lrBCAEtoItq8tLmXWYx+37+9tsENX2z+GgyOCZk90Z3A+PMJ
4MJrP4/S+XldHo4ZTJTCIumbuGjaypgMFnE9tiDfR/zSh5lc9p4ajXnnStLgo37Y
pJBsoU+Re9RpNeMY19buEBjciNd2XbQKH7qM/OeX7mrWieqJLeXiH+r3eEuy+CGs
rUn+ACRVfFEcI1dPPhfX5wQt56dG6BryoCml21MMdfh0Lk/8DUIoRsp7x6OI/DgP
QqJommeJKQ6Y6WzsTsQNgRjV/g3VhzXNFJotKbFtDoO40ho5DRAh9qxJHpblijeP
pjmTB4qtQ02bsd3StL/OUO2nmvGPNfPijlx3Zv8Ad1TvsJ850qm08kYdP7QgXP12
8ZfWtF4z4NBcWQLHlpqn7ikXwrmCS2gMXih6W+pWPCNSvuNrK7y6BJG4tMC2Zcz9
ojBG3dyp3SVrJRUCHRwnXH75n4+jb/lL+t7MJOje2u0s0Z8vPuTTX9Y/Lt2PrfUZ
L0BrSGaVS4AxA2w43V+rciWO9DBMf6o4sUzGQ7EAF0PNqXc/kNaB+1WjXoJK+QhU
kRAlqIQIxi99jp0StXopj+DU7S7IAJhrCGtOEX3YqB9MSjUnRsYD55um5p0Vs0Zb
usY4xjdqyEPCcjJib8yPl5np1kW2b8R32m6UJ+eIE9Kd4AkjqfRr+s44YVUTaCE1
Izm7CXWtlS10aaaywvl7iTsWGnCEs7FUmTlf9xdb3bHUYySPuhrbSKotalLFJERO
E/p4YLl6YN2VT2aMacUdSod0PoJB31hUV8JOhaFW3JPrFlii5JDTmeKRbAFrrO3T
x2HdmSVVyIDIoBGOJ2k7dAiyLvoTgCUo57jU61CcWkhVeo0RztVMUxN3TVy2B5DJ
LnjmWr+KA7IDi/dbbfS2Xte0NHP2qYgSfDyeKGIXbqkvA//R/0BISJcUWtucj8c6
0aA+2W2DIzWqczisP7NQQhfpvcVOMKOxaKaVKBrOdpnScQuZxg3gwW1fuTEyD1zj
MudUnRIT+gB7h/JrRjiW0ZcpmTZZhk3Miggh4CFs4RyI8ZT2PxNoOI1azpgkMBzQ
sLNQsdKqBvTOZw/A5CtdgoTTygf6zuv4SVSZV0JFUG00hwbMLtabrwP2YoXVJW2E
4oIV6+Q0xH4228oZSyPu80mdTHyJPdF0q0ug0dHz/OcrrS6pIBPSmehLGs+CTBoT
6rLIreoX5ZBVxZ2wQmNdKPCQAeqqLzzPq1jtP8XjKRdyYkAIMjvEDkkU5qVfOiGR
8NX6jc4eEYt0H0l889AYY+2BAFM+9DF2RY9rof7H4p1rcaejsZLXrzU4N7pEVC4l
Ek538fUK5DqR1faYV9sO/JnCz6mtwE4NSCSnHXrfe0WCvTdKSsdJh+0dsTvAIV7h
a0sHETb046oHv3WLrhOrhptUBNNRzdw8ie2GYDVfkA/zowL8h8PnfpXsiQGKEGhm
S5V5Qcc2cBuTFRluwZbIEVxsDOtJs0tl8nMchB4iG3SIJAj3RF0PaDhkBlW5BwR5
DaZH+s2wDFBZcj3ajmcanf6MtnEjhZy+mPn4LSQppwWK8xDt6Bcb48lHTJzihMyz
unrbDAn4CsLXzfTEpi+QdMkVzzy2jqx9MyGOW1lPGonrFpn/8Ohm4QAfLBSEqYPP
plnOKtnX30g0T5kqcPdsSdLT+Iht1ixw4PHOJRkpkHfD9e3cJsytkhoDJ8V0Kp6T
+rSfNOU/0oTnRAXJv2BM9+2llffA7Xl3uggNk24Q5LT5/j+d5oYBJI91/+2oot5e
LXfH+vmSTbuoQVRWITgWXX1CMmBr4I4MugtQZHNcd8qC1TKV5t/9jo3F3RLBk7Lj
QSokJldoYytxdb7HGhH3kIQ92KdIovD49+hej2LicGJRaw7Ut2A4kAGb4bpzpR6r
AVRhgWKUlNXiEum9k2ZGtt9lbghUSrRc+PVY0QuLSNbyBIbXeTFiZikfdXq6s0k/
g9lbN/Mvq9WbHu4/OrIOX6p+KH5Lt35DDM8Poex4QlQfCufAECAd2/XDP3FU/shA
SPbES6VvIZxLhrn7kh8+20Ur222H3hMo+3bB2rCIo+ddPnq0iMZA5Z375URqpHAL
gqFTQIBtIpSYDsumZp1H/8urr3pmdafSCTuUC60oxitbPNp8xWfnp5TabLDrsmpf
XcsFXB1/UPce2CigYpy06bmxQYvG4lXbeOfOX5B4Z/W7VjFxQNTIOBpEYSNHTn63
ayG5XcEKpG37FSEezqediZdo5BzGar87/Lg1eDtnmg+KMzB+zB0WC/wDW7JfAIoU
c6XyTBEBo6nwq/growdO0zcdE8zX4nvX0UqEU+JVFURjUbEDwgb86iAhTYzgQDLT
lcUAdVUDNpEAW7+5A1wqVO/4S0lNddAzDPjHA9SYaJiL/cYaxyRVvFF/sUzKxfPK
x5JpHa58TrTJK4slypRj3MEddQgzYGJrnL1OTuMpX4ZM2lHfS63JN3z/ls6s8UoN
8wJAsA4cfLPxAikPWK1wNHMKZSZjS2sHsOP56q3Fy9H/xYd2SCfTTHG1WcqA0XbD
om+qvtY5E8b99wnAkKq39hLa8JmQNiazEegjvV2Be5U159r6PMfLnizB1d163kya
cdHWRWS9tlc4xrUEK2/+78kaz5xE4dAnsCF98a+YuTvCAYeHDvJ0MK8j1XANuety
7prRI8v7yALXHxaKnr0MlY+TrTSzCvZzkvzOa8d1dcc9up5WKMjGB7Eub2dEXjWv
QoPz/79QSb/UdzuxdYT464NIvp7norVLMuqHt9tmuFCVhcjANsdYfYQYp/xsWtv/
DbLzRhXpk7lmB1yV7oIkEDyKwR/PmwJGFFeeYXWZVa7nEK25FDR+PFfb5c6CNRuC
lSydF5E2QLlYgs1Lfa3RPa80wBHcot9VHRVxppvQEyseA/b2tY1qJPa98dULiCJK
JN6nYhVVnkUkGyw6rXurR9UU5VUFwdgpbe4G4WwTnJbVMdj0wwT+btWZEoxktcQw
K+KoDRu1v8SrfOtOaDvKJjkts0F/3df5qAqj2HR5YE86TkR09g+Bnd5YXBtTwJaD
WzWo5jyMFiNUA6MlWKTDahAsLdFGHwI/iXklxZSPpNVXBagAUeKMLLFMjOnoK9RL
PCYj5MjcgOxBIZcng6H2ogAayjyCync9FRTvWwgbIwf2u0zdo6/DEwyL7iaj2Lkb
jfT4GVhAAPL/IHptyvQy7MDnexoaOz5o0KzMsV51rKrsKGDryXE1jFyKgcuu2ilZ
SkUxgc0Squb0BZ4dq3vfe3Skl6BjRdp50slJ3v8G22yKCjy1Zmi3B0JQnlgELY00
GZ4VmWNLNC8pu4B/PfwdZ9p0WHeZcRSBlsACl8iSoc1ULC6rLwdt3vT1uTK+Oip6
N2xyfd9nKTHD4hHunjivXnCxY1o20M9IGm+asXmzfqO9ODzQCSsL4JpctYE+qbkV
qRwgOgVENrLIGilzfvdhN8I89eZ+xxPpYhgH2/hU7F2d0CY6vyzNHDyoWsHJBcoi
4keI/USczix7BBJblP6g3Bceg7yJKtAedt4+ZB1mfL2y+Ksj8vAudSy2Ar0tu3uD
kdsdHp5K5lRw6T+xIExYUuENPDG/A8rSQnq6tA1rssvbimQWGNgoLH3jRLo3DQXg
HX/K8RYAIwpmuhWJuwPosgtxAD1wMVdSUzyI8FZkGYgSnsK8ghxXqlqvdK6MBOQn
F4d4Kw4nG3ul0HtQrvgOqktD2BapazOHHWlouKPPO11rb6AYGWOGgynJgq6uAp6d
Lp76tSBZqPOEHc4qNd6oq15k8y0U4wLferwZjtxxCQxL3T08TyunMEa2L93CIbUQ
XFI2dtBVj0L4681OqEg99QXDSarDz8MRTAgww4ysEpGyXpYOSbBsICX0TKRgFwBo
KKc7eobbLxi1Mh2vFiWAQ/JKuEIoCcei9Wuk8M1BpoxngLeklzNhSJ0qOsP5exxh
pDRiyKaw+MfkAM89VW3K4eTL/Idf9xXxHtsfeHAN/aXb9lS1y7lBBNUyjKxuxg+Y
wNv5ALl2vgbm1zglycgAlKYNAmHVr7zBwkNtHm0piXzyyF4D+uQxFTk0E1yHCG4H
1emAnjT/NiV16QIngBRWssDUatQfIeweM/6RFkcy05fB9YjUZ2qhxfIT6ZphAAcu
tToa4w7XySe90pq+S+iRkG/V2J5hi4eSud67dd6Mwp2drlnjeNo0EHssYDl6ic9n
BCtI9259PfxPDaF0+3JM4VjpiFIEip+dxkEWOx0A2IhsjYKbZYT12yW9GHsXQaJT
av51eNqGaxm6PDrfO6px84CqfbJIvfA+cI2ozEHSSlefXVqMEuvPhU0eJNlbwWr1
AjuswLzheweT041Xv8NPOP9N+3Q0hjPgHFAx9Cb9Nnnkh1EisjbXZEGTo5mWZkeI
AstNtukI7HKkdVpHfKePRPI51G9OQrYnybilBCyGfPBkR+QWer+knBtLWO0bflPZ
PZ6v+W6I7ngTpApSmKuzJuLQwYPM3J0O3oi2594o08L/5PEdrEz3IZPhk99/CMKC
cpDI+53HDkDkyt8kJg9yJ5W7Z75L9FK/f4iSPnL1SnbCKFxzOsaNBI3VNwGDKIsm
YBsbF6I5f7Q0YB9RC3b5dBUFSXKe1H6iy7tAvvFJPFCGTcOTFa529Pg8vwJhAxXX
LAzNoZqosvpkqwqDtEfx6JmE81+5tMxzV4NTSBw8mJhQhLZ1Deeg9RxeWlekoO+1
rKVaXowCeawzCfiikPcQq9d4DLfV9szLbJOvjA1QyE4BXLTE+Z2ascLuXXIG1Xeb
/ODYfihj2cjIlAmqf57kR7yY2d9ukAzk0RdbGatN0PpFFd4vEv50RKGSWZ0d77u9
vwULrm4B8nDvuyUJuNd/VbT7y8oOkfjHp6BmVdeCQN7dbTVoQeYZKgnP1wR0wbC1
R1dd74MAorP1yh4ocfM2jvd6Rl4eq0ljE2uxR1f/zIXu3kKa5aDIKRKXdWD7DX8Y
hfdon2vWZJHrKl/qf29vISGBczhKRJk/wzUxl3RhqSzStA5otC3vmovQs2W725j4
LqgbdqOzJq2KEclWlY/GmyAcQE15dZJxIg+gBhZMu1tjNkJGEgm8SjqqzxbRgfwE
FqneO/VlfhMh9+OKGWZeVSQqgCIgEXBA0+WSWiY0tLK69gKAICoCNKW1SOf4fUXU
A84Nd7xIGzE4h11F1g+FmNtNR1VBC5cvNaaj6Pclss38o80JVzjY9Nm0HpphCX+W
32dI0Z8K2ER5avQR1qbYH6hV+enAy2KsnjL26pXjJjFUKemL9RV5p+kSFfj6w0tO
oM1/fBaQWsQao3ybDepJQp4cxFTDYbAhcyUG88QDfdMtPjfEwqTVZXhgQ+6Q031b
5T5GlYbi+eSxEq/n8PfIjoLbRyln2sdG8jrCjxfUNcCGXwU00C6nrYJJKVgZPgw2
nBlE/yTtlHHynuq759T0nioBgYwRZINy08LpXjPUwKnAQUfLtKNsEAVP+9nzVwk7
Y9p4d/agksGp79jK94CAjMwRA3tLKabwQX+jnkgfs/3RTtt8SlrPWjNmWlAT+D0w
nrlOucreLcblfYzgVJwP2OEv8R1U0qa/d4LzNhrDWy3eMDMLL/gCUbGkClVF9YPQ
6AONOVExyvwCJz4SFjNRPmllvdmoaplaC2c4OYAvftkUFqx4cBwFXH5bsm/+opNZ
zy9tTxBGYY7J6s36tQwnOsHd5ZsOsEBuWcvTVeTBzcAuFXE+A4kiQVR5SlMejx8S
IRf/hwVvJG+qSfGQ5gNOG7LownSVPggPk/KFPyMr7xZNBV/fjIRVF8vk4fo1uFG4
wG08wGJw7fp+tPwzHVuVZ2IDf4XPZkj75196115stJZnudVKTS1FUfZ8lE86ON33
UxMyX4xFPnn7Z+FeK6pijnPV+rPXdVLOVnL9OafOj7MoSO7A+Kp116IrmRW4iycZ
3rLyybru2LhhWmy8h1vZTxj/s7AWx8WXtms6g+dqGslgzFyfuS7olqYIB6mxJX8M
HANsI0mqdJs5jImoa/3foEPhvwYigDbQwGPJRTAzQwCcn4JV0sw7dkjn2rtM8VDq
k10HnfDx1wZojYaq21pO3f/t3YOze4aos6r29WOJrx43W9P2mpAhKODFNKQVeugL
SyLPJKHH4mnDmAaaBT1bIqQwudY+GQXKLA+ruslfscGY0DRiZMzHyFWsHEDKH0xo
+nSkjblYKtIeUtXyov8Dz1FrESX2oJAVhZk6q5X3yVHTn3EgnZxrs6V2kaiA707A
r6qsuXkhc9Rw/DH670na8wWoaQjhBtDxYZZ0NSinAJJee/EvBuiI7QdduN0Gt6mR
ensz5eyeIAXHmQMoC4unYZI2Aiv4/XLkn0c/sUdilESwx9v2MGe8egLF+U3WTkqY
Grki5a+LCrDFR0BhMJ1i/Ey3yntwP3aCDs+0rzj7VU9WVHFd7PpeTCbT7KdLm3wY
kn0rj29iv3DL3lgAs52+84nYBejxM0XoLYHkTl6emeQgSU6mrklfb/At27Nbqprw
844ekm2XGLKKo/BAe9mAIwccVYR2RWjSK43iR79wf3LNjAyqhWZ94bKBiA7AoCnc
YodJ5pKYbOWNKRipx03vjJP2CuE4zke3gfgEYZIlZ7xPHmXU67zJ5cobu19Ajzlr
sDhI2T9OcCISKKjz+hj/CKf9kdkr2rMyYLkr8WotnKaLUwBA+uBRh2iVeNS72YdA
nNLrQ3bf3XPu78Y/WEHB+n7x+XSnxTwiKo3xQroXkrPu2TsQvng85h3bBzvWfUtF
+tNY+mLDbW69VJwrXgwb14LJU7YPT3qmWW0XB0AU2QQoFxI8X3qWFiojkzJIA0Oy
deaWMcTbx/JH83JsAbf8giz0kP7DIH6ST3judyi5i5/89aSwavTSdXk2j/BG6/Ig
cBCMW3W1obo10wL921tNCg9fPngMtmvWSLpns009JQBexE5WAJxh+H1zb41g+drm
bOQjWBuV3XCbY6l1l08QuPnsQgsR1vsaf93OrUEqAB2CiSPPcgR6CLBxMtm3GBqt
VdBvcUcBzlbTNOPXIF+TOjBZC0GndORh+8QoMNoGS4nZtmBTsCrtNx1w7FoY0y+u
CWOqwoJMj+ssRPpsuAjaBKppZEpwltaRPJaK/V1MZ27O7NFQYqAoxpiWjCcz3nFg
uZ3S6YV0NAr2+d+3WbMY665kRgaUPRw9KduqPWwLKlQcp5381tu9hTj2do7ReFOk
HcavXcQnezeC2Wz+DKhxTVJEV6lpvD53dahqkEtF9/6k4XV5OhbFabXnzhFM4/Ia
RB2OCx0oxrBLFhOTYW7QnqENj6ue1ofA9A6W4XMhM2z5Fu0IPg2vUXmoax4Ordmp
M5PinGCN/09vKa7uOol1CHz5LJRi/tmU+SQiEEkw2+C2aMiL9s6Hekb4ux7HyVdZ
TgxNieB1OUYm8lFANU3wsAyDIzbNaNJ6y+LIqwMug4LiPaEcJeAWTJ5VquhO7Cxw
TbK2QvwvHDCGnghR1rHA+eZg+da4DQxL5cVdR/t6sMN9wehL5sqU9BHFzB8JhBSV
IgNEyUqBWPQW0M1HHLJr9EKJpxNgER38m8Tgike7JDv4E1fxqMCDBFKFuKdVJwzk
lSnZ0ehItQbniXBaUICQcIwv54oWjUgkSQVmT9jStSlhllFSHIToQ5RihFpxK337
EXs5g0A6KwZeg7rabHgtbMo74ziqBsRHdq9ee88r5mAyVjKHWgvyJTOyj9ZoEvRd
cyv36nKeIG45xOnsKs8E4z0xD2wvxd+Uy0nKyKbu6yfsZrIlLWpOu3fUyzfb5s4k
HPydFZFSBFaIvhFVtCn85g5bhmlDJPtwUCVAUcT85f+cpmJKv8pFYb+EuvcNb2BX
EC4To4RTuGpgsSS5pcE0qG9ArBCT1ZGhZf+YnaugLnFgvQVqgOwpFe1hIhNYiYOY
gw4DsFhWrFAWgw81Emi2SCy62nW/c0IcRmw6auuA2aeiCHBALjF4Dy5kwK2O/Qio
ZnhmkJITynUtBb2671spdmMr6UzhByk6US/NUBOJuNClsRQYCkTzLibJAGWUiGSx
z+I9l/H0KTa1BSU9McYktATedyTxC/syAPAIsSvL26QLgz2QiQ2lWA77uvsSmk/j
lR+/g2zTDXKaB6+PsP2Uk+RrBxe6GcvUbHCQT2XFn6/QgEN3Z/JDbx+1UWo5F/sZ
01AJIxZQLJ++aJmjkwHLeLuFFnXTi8sLTEYxS5U0GFHcm6lg21MLKfJBSa+Yi2HE
Lv4IhBdpWUpLrJQV+ul3mZqZRNXozK1U9tQjzHOhoI50iXJxgExsT178SfLhCCTp
a+U9K0jxSUOsYoaCj36gdbRmmfJ5hTGf/XvCOwDqVYOYkYTccDybUpuh91LSP4zA
huEnU3rRXGrCi0cp+zePzPLv3ZxwYFY2MHpv36EX0l0sYU2W6OgY3MT2iGUam1dH
+b7VZYYqf5E1wP7nkIVEya8emmHVveFGuBFCamhg4aDqj5CnPN6QYYjBCf2IhZ1x
OAjMVEqgJNlovOnef6lsjvEoktrbrfS9NtJQoV1eX6FL5kzINHzkUQg3KphHQT20
5u30DkwqYy+n3T/siCBnyTiBoRVGqO0276xxw7laDjNEB35X45jncK67Frxic+Vy
jh1exRCTROHEBU/N3/uejr2t0g5qsibUo6/wL6xCo2GVDK84JjeT/hMf0vyRVP7U
LdEfXziHvg32KFULt0FD7h6tNTE9hsUZUGg615uwbvAdnRaTftMamkqDJSjFGxqs
IvSzrzh7w3SlMVYONXIqwQCbya+Sdw6woKckXv97dC/2gvB3xbqS/grlpVmNhl0q
lPDEcDMVAORYG8fgsYvPqyxnH7MFvWi2Gd32aVAckZ+gcwOg/ZBL8b/y2EN/Jze9
uMAxFD8IkrigmKn2abUD3wKiZ/DbhP7Q4qMpQ8EImDLkoWz1wC/VlFlDnXqM1StY
mR2cyxBuLOklguMnBq+2FYKoPojOy8BG3n8U0nz4gQmhmBeuNCL3Hjl8g+BejiY+
CEkvGXJgEYM8IUbxGn6G7sOCu9jGtjEwPVqowIc5Ehww6Mn1XpczfKroTxC6PEsZ
kilX6Yh61OV6Mi+OplemUMZO+7qSB5tRvylSOFG/RGkw1vV+3+lwC2/cx3rEy6sE
EaE46pQTpLiDrC15Y7fxNkO1VrnoqrDNoF6pOs/g5wwSppC9zsvo3yRxgLxPFgai
UzzK89+m+WuVYeyt58WtbJ4ZUdsGCZ4b32T8Ecw6JutXUXmwd6WvSPLj7c5DaTTd
IK4ToLuEkTJYz4E5RilItop8vGb/wRaSEKMcmcKS5lnRkUX3vAFaKS8fQJG7b5Rc
wS+LLIrOYpnzGIusMzfAcQGXW3cMeeG2BMBAiGXmE9SA/VhniMaFQky+IK/4jf0j
gEI7VAfw9OwFQB50Sl0mhe1zvzTofOPyRr/0Y1cxUhwsuXgwZrPC7HgYypjQnL8x
Me/lSAnoFvLFqZAZD+JTt16ecdNMB2Zx86E4k+vIMEx4wmtDPZtaz/gVWgOs3pPK
MHZPdDTCBFYH+ZBqyXJnmUt4WgBdLbpKqiYI1CyQEQC3IJCb2ePpAZ232NnNh2EV
joogtWjlP1lbr6sLUC/FG9Tp5u9Qd+cDesMY/hXmLKA8lXRQTRq+ppjRqpeNXNe8
Ez9FkTiijj1eI7UNB923fW1ksnJJcVi+/ORMAftAZN2DIPJKj8vNfvu+cqFi8hw/
2LGKA0d7wmZhc+qKJGDaIYJsP7wEmpWIr25TXNMBUGuxE2ahw1uncZUlNQeqDiWE
PBfUAS81gSCiUgumgimUgDKuZimuWb229EizhYvSYUN/QFOgQfFf8KNzTrqW7Yct
QTZfkPFpe81/Up64L+KhPV4lrAlVqoCtd8q+ttNa8TyfeC+MYPZJM+1qYBsRcW49
WWzgo69C+yAOSl/lWfzsGcDhiAUCOp5XsqzD5cuxI4qwh0V8CfW7uUYFA8vPGjaw
DujVHRStZDvovOmQuDh5Weg5l46obA+Q6pN1LnS3ZvqWsijKToCZRZ0VOqNn0bAU
+EEqgCowMHLL6Mot0N1qRpCuFWEPvKukSamdmAu3FejWp0cIzr+Qt/jan7m1zTSB
3SqBmJB0udIl3z4jNz5uz2IfYLQVP0DBR9FyLSMS1DiG1SgjnplTKVBJF0Ny9tMw
l5L1hfXzP7+OB8ERWll+kKIvvE0pGPo+Pmsc6AXZpJmTGo2zk2yMj2Xv2DAW6sw2
UZc4ZVfPFO5K2Vs8WRXphTs3cpO6Dc/gqYD467UTst/oCvHFHnelVS7Mgw6PCRin
FVZBncJjZ63/9MESxQVS1e5wxefONaFCCMVW9gCRQCe3QmrOL/Cq2pZms5YV0p1p
qOl1mjeAM30xSEk3ooeB3EbGPC3aj5bxY3wvO7sFURQ0tF7oOSpwMfyXH4ai7nQk
P0Z2JF+l4P6lEYg7Hs3LsAbA5E9IVvh90/XD+X9+C4fr8Q1Ekg8dEU+mLk87ECKB
slqrkBUdk4TxvnIEdPRpC+44HoFED3puBx4h+AFKcwaf9i7YV7vUEhAjkOCF+B2Q
Ld0WcGG1E/FEcZ4nVuyfZA+6KgGB9F1raWbtiZpwTHLhLdNXvFjMzm51OOzxduAy
ql6OztawehE0rcVcxQSEmRWLmc+yVn5aeY8CN8+aBRuswsFyloEth0++7Y7C9LEc
W0QhQeCCtk0Z9YNkWyH6dIhHzACici5v8zwoXzkDyC5QDbvJo8rINMHd0o/ZOMbM
1nJXuyCRoWFohVuvWESiaR75YDVG7DSmEImAac1lOUVt99GRRtXCNMJj4KTFDudM
QdD/1wjEN/2phPMIHQ+nv7cSxC0pxA65AfXGbEv/TLxdC81Pt8/DnIAfMHzHcEap
ZrkQVctcJwYG+9svymtCTcXcNRfXn58d6beKIZfX1blnH0ydQtwxHNOaiKcUJzUt
saRmkdKDRHKzhGtmc9dF8heAGg5fcyWwMmVc3cpvrvshMKO8oI1I7RKTZotOj9xP
gKXcmDo5QQCyqHcbADUlThostRkWzbRlAKkt/iZA0++X7FOHRjnV3ZPd90iG/9MU
LFTdRXpDJzCmeKdeEXavgDKfUji7I1ojQVIysW8hfZcr0W7sGZAYKYljag3YMu2s
Uu0DgJ/WZj6PaV2DhOJ3oMSHf8E+chjgThZCOOdYKoWGunRwxGV4VjD29v2PvG9l
dVTlzXX8PO0iR5awWogH7figEmwH+7mG/4PRdx+pc9F3fAtGmjvHZRdD4tx9/HEl
ZovCctrMJOmLJe13CVJC3/b0shz994azGz5a/ysGFck/jJo2BDYGWJTL/aZe4kmO
0Kf9uCjJu4PEZPgLylXTNx4ff2Z9Z6HT4nxs1fV2TE4ex9SLn3AGTKsKjC1XIR6W
v3P3awqiFbYV2l0w+PfgQDPOxLeZn8qKzm5/OhY970fUNs73tNKG5/ChWfyc5b0y
KJYDRKdSbCcuik0qvr7Myk8JYQn5HqcTD+o2Tme6moq3NOdkm9PFDOmAXV2MqN3k
+2xJ7JFv5xy3jdZ0PPZayB+yS94iLoQgSA9Jh1jv/IDVgR7YPiNBo5FKJzlX1fxZ
fn05/f4lBBws2CPfyBz+girqtM5rHkMVPGWmMoKaBfV+n+3cCKZ3CqefrSYIhd4+
jyt5lQFvZYi2p0zZnpIOSxN0srzqjo7hJSLYBS2Y5UaKUiyjDxWhiJj/HSWK/Pef
GUZmeKUFJCA4QuFggQ7jm0Dy0so+87TtkhLBg4si9PyINiThwWruXQ1haaMBX6G1
J7g2T2H4m1Zt+QHWUiUPIoq8fySvmMsc4MXDT3r3+LIfdRDdAPy3iSlMs7/oCW9u
M8uBXgpeTrQAl/VS3qYjSGC/NNd7FkFB5cguG5G7Jol7LE6KutZh/BST/1h3tKV2
KbFITZM8eLS3ONdGom+R/PqZKKXddsGuoa8erX8PDaZ5c5t6wGEsvlibArc7bD8W
rMwitaXSXtCbk0z/8RxaYOQ3I2G8aqMkoYPyObCd5jUDVFJXd4vTMIEMKbY3RKEB
h3KJFy1z7wf0LIxWFARgsLGyErBWqq9oRFEDQZz5C+3GSeR1xsq0mhB5vhleZOs1
nNn+rtpRfmCUtguzXlLK6IxbZiQ/jEHJ9w9vjUjSa+DhNWZSBTt9zGOqZJ7Wy7oh
nHLe+HihHbVUm5t+ss/TS4v+Wj1iwiLrwaioFGz2aI79z4d1b0AIroywQs/QVMCT
61Pc0vQSa0SZT3tfA/G29kkIJNBt9Kr2MmGO8VCkLSUuu9j5AWGhLanvI6OUMu0P
q44RW31toc8DoTOWV2DUYpRqi9xqSyI8+tEZXbAgycuLk/kPo65wZDxBYqURHf33
ty+1ulgEsNRQAkIn7FL0RDk+kiEHte3rU1mVh41hz7ons95j/pJCow4fIKMXWV9U
e6Gw3TmQX7fDvNBDho/OvfySQ5WrzxzzuLUtGhlw/kITEB5BwlcFDGASAd07cPTR
T8d8+vRJu8hWnUcWx3wMbZCnPoRxQBSeV61inVXH7Y7GpIoi3KoF+VBi39JV6x4W
9VYbUQevWNYeLociWFhxr1ylOxryNlaiiv8Y3oF+tAI7XwNEr/SUDFVEYuXjX2kC
cakw3O1pKwa9r5gGUpTxlvm0xgCJQr412cOOlMNkDjDuzfflDZ28C+dKv0MqFwaP
0xMFHAPR/sKIAFXEG1nDwqVdimkGiuiFcybCYsPsqjJpoRl7UdJg5vUGayqZMxhb
Qy8HoErk2Py+d99Zj32vcHcV8EOSOnjgAqQPRX9Jr4uNv1Fq0Nh76skG5Ghn92wv
immQepLlN+te61ceA0kIhH3Ftacfa+cvkYYdRcIbRwnnYwoe1OGePt6M7gYGd0sl
eOrdrgfpDem/BB9oweFxloiTUeLwqOJ6m4De5lGCFk8gTzD2jrwVqHSCvoMGTOCB
nQZ0I5J+x8bosnrRwI1FMheFoKwQQAUwuoERSscB7B+oG7ffmj3yy4XSaXRAI2kS
b+Qehx+a9IACCEHXz1jdju7CWdRbVcdn01xB0J5HufHR/EZPBSejZC7ShOCrsiaU
YxRA+IOOQPn9/3JImvsi9iiNWhls5LzQ2aRAXL5Gicb2hp3Y5vrv8sOcs7fxP7HS
hmwq1rv3v+SejY1rq4OPMoc4EmsogqKYro4uvrJjoAkZbdqd2Ma8YwUw15ZaaYUM
qoFYcFSr5STMFt5Y/XZ02LJPwOYNwwDL2pqAQoiAPKAMuyVZs5NMSrLLmyhmRlS7
lV7nsybVVX0m1+XGwq1JvAhwI2YLuqPYrWwLY4yzAHUCJwihkQQZyImx62nJW+Tz
zhbQbnWWyyekqpNorLtwzR4kRBVirWNONWT2WxtZ415HyUXYZ6cKoLIjWiJLdtBv
RC01azsT2e+pKmZRVgonKk3V8hwdGWJ2U/73HGjJCyTmTsRh3iN/0zLaCLULjvwL
IRmWbKF50XDlzTrzgzb/td/hWXe/5k7yecf57NDbY+PH55qnf3/zkCIfwRoMNjek
Q7kSaDK925l2aQwwCOtYC/JPsQw4dlRtclijpiqxWmSjn6+qra2R55UpPlsZMFc9
AS3TIpGCVmEOQwxqdNjB02Ba9U6A8+Pn2lsIPxG2khFJbhOHWBL5aBsrVNvp+/cG
MLEU88kBMx7Oj8hkEYR8iyokJHlQcCBSARD9ScOUq/aHqxAHX3TMDfcB2Fs35P1g
4/ylhsM/QDnrkJyMxanmG7C0yYg4AfC1f8Rk3YkiT725PQvLc5yN7kMwyGqTOmGv
ZGS/SedOVzenw2Epyjh5sq5R1M1WnjvrQp/PlY9w2bNh6gBkrRfkihgLAaxOYq5f
PLDu3kpz677+4kmEDYcYlHP3QUI3Ki1oKIhm4stbO9u4CGh4arlyf1yiztIazyWc
4vo5HwEVjIgDWNeocOJqQep68oaZ6g1u5qk8/fXsNfPdUl5aX3hbjRWOIJOGHfMU
hp+5k+F1xXXGzBs5BKUy1h0f3yZfIdDPsO3aFjbdRWL4YAWh8kDmQfhTJbRIYFva
v/qPUcje7SmFtzHLiiTu3yPgLpxkW1WdvLfdNBiTpuUZ1geG1/dqMxVjQ/0un625
1+FkGXJ6zVmzdqIUCxx7MOGGPsH1EsVpvmXHtIWgtSIb07Km/AHkGKD2ntd1cijJ
tnfDN8XWkt/V2I9k3YwcIxCWSQqp/YcrGOJGZEMdvc42DC2sebhB25P/p9tuzQeX
/rPqi9sRPiLQe1OLOWAg8cvXeHgMuhmBLhlLp+aD+HqCI/4emMtSf83eECqC18Ce
oKgPQbF1zf6FPcKi8AJXYzSrJ0j8Sebz4Npu/o9teXc6VrMyRaNAjVJN4N+Pp2ez
EfcbrVsLmLjao24xvABDg4uiq817NHq/keaKiSWQdb5mgfyDtg8rZqf/eRY22ouk
qdYXg+6qdga+SEJUQBz0UnnLWVqr7F4MXN0om2qKpI70pAxVFIZnkowEYjpDb/DL
yhf2mlyOfcQtZv5JtzT6TuryonJ5D1rs/qt+8q6EF5iTZOao2ALf4s9RGkj2q3JH
p8YWS4HcwKoUS39ed+wWDkxM5XdFAZyuuoC1poRchsC+A9c7LBIJbogiENYyoo0P
ZptU471s+f8eZ+Lyq968hixMsBdtX0Vvp39XslsThgq3Rn8kC4ImFP/Jw0cEmUQ1
hZmWYCRpOtPjzY+mKA98ftH6aB+ClI6SbcujlTpTPIbLv9eTgkJNl37GRnuYxjGe
mqGMM9iCituYeyJzFg4zzn3GV1TueX03dSA4IGLavl6YWHu7v/7TSaJ4/+CeWt0P
BJFfmSDSKSywlLfVC7xLSKE8SQegFGoXoazuXX8+GCXYVfhBAxe7ooBMTbYKos8d
Vz2SpyPDsw2wWLaZYnAWCITqtYluwx1m8B65uBgCIUP4HqQetKl95hY7A5kx8ysm
M/VDBgrE7dYhTkIDMftj1PYIl7oFAbOw8GjSKPal32daPFXeWZKKwtiCRIAYuZUd
THj7+/GMKdN9F7kj1v9yXw6ITwqOLNoyoJ9oiyuw+RY57AGuUbYH9pCdp4jjVtyY
txbG8bcrYHz1SNYzIutX27l/Tp15IWuAsrccGxcHGcm51zJJPVcNZkZYKslRvULN
XW7Z5xSpkJwD3Q+kY1/xHoI8wsjS9R0sydlAS2d96xlRFpPMH1YEiaebmqgNmJET
YNDYp93YvBnuh51I0/F650jZGqULwq/ND8iTgkpdhJ9L09KLdJiakcXR9E9AqVu1
yziDCFXvA2nkCnusRP78fqKgake531PIXH1hJEpvwms3wnWr39oeSqBk7nn6xVor
2YZoXlMe7MEAxt2PZKRiV8a1B/C8Y1rENLLkjDB4FjOSy1ICv4h6usZf7x4C4RM/
HAh0UMr7N2XDIVbwesw/taoCNlQZO96ObIFMI9BFRzyQjTyRPRN6OvAYDO008kd9
uKoZalbPGRt8sWeziOEiO0OQiA476Lu4Nvsu+4XAGPat6d60vOI9J5E7dWjcPt1y
Il+bzBjZ5GmHaFEnSwcRD7+LUtQr83FvGubbRl7bRApQTh44xrjHpCB7Z7Q1UB5i
f1riiYmAHS+ei0ww4TvMmXoA9jTfWz3Kv+V8C+lIqMAXq8mUSeRHkitIFEjunlUM
BDcnKcZT0UVSlXmXCwUpeEPsG2CuMjJiC48HSVrX4EDkegEzXmL/2AA8yu+t+cHd
VC8nNQoG+wg2C1s++2t8z742+40wrFvTzllGShw/ilFE/MRF0uHAt1xbmPa/Fc4H
q0Hzrtjbdiunds99NAYAHaFTcOWgAkHaD/lgUKfLKpfH+k5AQvQUyccJgHtdNzA2
XY9CWe/bIheVd5/PBcxoXeiLiU2YfOnFAwLy71PPAWL4MaaT2vMGjfdhz3aZa27w
Kbo89o+Re95r2juGJy8PjPtRApdrWPsWnEM/H2mfOr6nkse0n0glfAXkd0pR68oX
jyUjC5lD6qpJDdV9VLQ+/uVYXCKCLxleM2CcxmuP1W+eh6R7AWK+MDhTEe1IWZvZ
Qzo8W65+/7MF4YbjjQtHg2IHa2WDo+sl3Ywev5JFEcRd68ZaIpoJyZb7qkl/4Vq/
Y2jkSrQdP8kAMAcO6jCQCDfcmIVWp762wG44VfwjlsJzaHJ3KGQaF6RHFt4oG+M+
23LQgq9TXLllBRS7b3+nUJCr2eAPE0b3LgPboq3ErWr24fdPnRmz7G0m4u8HaCUo
S3JqrLeuNUK2SuLcSZ0Llq96Yg9qbbft0tfZ7MJ/Wyrc01eEmMigPh3s48itLjZ6
0F81IFVxOU+TnMEG+gQR7ecCV+Pa6HN98YXD3XxSCqKFo9TX9W/8KNDgzy5SxLpX
RIDrGg0E93YjoJ8/RFEBcPH/JW2mgT5dbU8W+IBsE3WJ+76Et1ekHfiwXaBZRVkq
TpebA4P+IOU90pj2bH+FWPTpuMA7VFv2NmqmxVjlPLkZJVdXi6G59JTeUebLqHFl
BTgnE+ZqSy4rVy1896jTOq6twdKF8FB9braFAkSHBVMA+IKIOH7R6nSqUZ7ywU+Y
hs0ksRr7nF1d/F9x94I/4qKrUX5hdnH3asfOjKip0EJwcHavxY1BNKlvgM/zBn/p
+V6pE9JDwRkPsLxp6oNouFX/1p/wiANu6KC4PZwCyB+ejmxB1x9oERr2xJiOFqhG
dz6hC6D7/x0arToeEmWXymuY7Et4tThErtPse/aAEQYqC9kbtBG4cj95cqqvBH+q
H1RkyYEfPsPScflsW+6jy03kGHWvx6AJg+NbgnU5So53WVd82h1P/RGqQ0A98G6r
Xbmbxtr+s5suS2CkEa4FCJGQJMnFhACXTPCltKzWq7kI+5euJSds67Uhjt+iQG0X
uxR8lg4BEwM4YNVZUmzhd4vHsqVVTzubCwNWJ7zitb967ZM4BqAGWKN1cUFvRorA
9yKPRj+twsckn3XhcSLJsZ2Oj8NDCePdtfoOC6RrNLy/JnpoOQQCvU1BGwR8XhST
eJuG1okGaxeaTY0XXXkoum6JsEsF4jOK5f1/PrSvCOw9TSw1LF6Kkm067Q4j3BXG
u+ngh3ki+VoPMiu8lwBR9VPcCrGLV3+pln30HQyPLAlvJQ7FsAQYA5J0Vsws825i
uE7PH6mZy8lgmmJjxTCq3w+aMYyNM3UeLSGKZmFgvsm2UVguoA3DUjvEq929vD18
diRYsd4nCEra9EUjeWhgYbINc2R3Uki/gOlQtCZcoK9EZrJWYqeE2Vh1xxER4ApD
5rKPPVVsgi62NqRnXynlChMoVBuAFDRNwV252qfwzSGiIAgTBxUgubcFFqs5kH7J
UKN4yb3tZQl/lb2wDWUej6m0KeIJiptqH/ByJevisQweTeALlS2u/bt2sBzg+Jgv
maDnqC6TKtfMJo6T0bEMur9hxbHeUF+HF9fSBSsqgJudXCcj2VRHDW3LiUnnH61J
PAm33lQEb7N8714Rq9q0Zwby1NdGfMO73V9tWXL+0pqdjuuaCzIzM/gSWzxOzWpu
EpB95BODcoJkAhnbDx5j75qqMjbJCvJ24GrgUx+V1rdsftrpqaQuD13TBHLC3Ixj
HEVvhVPzF1kI0u3rrKW4N+XAmRFx/CM9epp9RMaZniLSw2+MVdurg49h6ppsqrIu
R8mMWGyK5QYj7aTnNQXsy+Bt/E+6y7YCkrIcGEshBi2apKVfBktus2BKbG/37SjM
3MoF3QMVGZMZmZ7+GKQcSxIkeoyYeC+V+Z/fUjkjdEtcw2LIWjwhHCtaoEQNfSDZ
+E1h5LK0Dw/8lgtZ7gIyCpx3Zb2UvYYKR0Xc2sth7yv+XUdxUJsZFB5EuaSjUUMd
eXa1m0Z27XcrS2iwHfFa0dHRHdzudxn3ySGklLNH3LWIaD+cc1bNmdMtc5FNnzxa
9xbD0G9ZKUA3ZUVx0+vtEf4uCYsp7PVCcvVze6lAJV6BN9tzvZRJcKHssTtswBCW
fsgGw5WGmcqhzzIQdPJhJXokceDSjFek9mfd4QY/v9h9mu7iPomjjqfV3d9fW16b
P2e6LLZZYIRr76Kie9FdZl/noLsg+7cm2Lz3VJHT1C8iFJMqt8zzIq8pDnldASD8
1Ff0G9rVmgyDIyTmN3l9QGcUK9BscRB7JUU4qSzByWraOCOddzlLGh4diHrDWXHe
jZFKQs1jEPK8SpdlEAn8zblvRovRCkjUBEfL3S6XmuOtBp6yOQ3q/SLxp+fJPGGr
6NsKWFCVR5eKsDi7yN53lls9Ge8ihpWSZ+Ddh7Q/G2AhCN9AitIfx4fCxR+ui3yr
QiRm2aEq7ZvMm2sYcVc7aRZxEOc2JXv8LAUVJmoIC5IsF4H3HnmMp3qGx4w2xHrG
Uu52XJ3Qzf1Zb5+9oh79KKpFDkAk9F6XyXDkXpYMb0MsNiwfql57XC9AsPXR+Une
j6lD6fpTIm3L4++CtpphPkEvwM5tSLzQc/Jiqr6oSWgk/Ua4P8QzbKIASOiZkSHQ
AOO8pJr8YDA0JWtt42koYf4qFVQV0N7q801+0fRuUTEevDx8utrk1Kp9y1IVjA4D
kIiGsT2wbMniuaPAlff9txM3wFgTQRg40aBbcglLi6PAbpgLXZwXTCbx2mfUGZrq
E/nnw/cYO8RWkHf827VTR3sL7ZeY1P+Fu20j4umfS8l28RG/39bq6fElfGWNNvII
wVQ9po0JT9iWxBoQhGBXhO9ybp72BEh6/A9GMfgCsSOh39V0AT+ldGTC5R4zXe5L
mMKwwH7uo2G08lVaACl7UiObRFDKctQkZDzNH1C5b/6N3QCcrACwGyRtGOdWLz+4
cx941RgYnLkpuMGpWiHyZE1kYMZvnsgR+oaPVB187Mlu6VsyPcR6Tf8uv0K2AXw6
v77/5Z4dY0zQqyIZFHz0ORI0Xz8ox2cCqOiQ0afrW6t9zfaO5G/BXAYwhgmBOQYk
0xX9cE5IzqyJ1iTtsRQxKCrQiB+joX2FD/kKqJMIH/9mFxLyD5EvLm5zqJ7siwIo
VFH9qRadT9EDhUsMXda4jehgwCQxDfUSc4I7XjM69GN1KevkCjbPrLhF2JRSFclF
9VRoWwYA5eBwdVm1eJiHD1ih6KzfBhETU3HT9HLxj9fIhDZlTAjD4x5du/Podwpt
ZYwrhlatovYQ4/3o8HqWvGcZLsb8ECNJxbE+XQTksvwnSa0ZYbOYegGwQqKXYlgn
lMdp1kP98lIVsfBh3nk6tHXJhG8exmkrvZ97fEHrMjuh2lVS1BgAOCzT5jyCd3f7
iY78uSyG/g5/QHO7bVgGmraQ71IGPDS1yThRHVNLHWJ4CxS54w+r2lcGzbyOQ79K
ncn8BLc2sKigjxifVq0Ksn9L8l4f0JQhnyxO/VdUVRJFaP6pTJM9jNPRHFxlRldx
QhD9U5nuFtHLh8XfeTTaZYms1olM16uMJ4LyXdN8lfuNmgLaQFocN9TlNgY8rn7I
mBlxLJQdAo+dNtEZJ/8D+PzMIM3WnsQia8ybCXhyk0MkinthIb5ZleFMyO7YWUVo
xcC/kzRCUqPCpS3hmsKDe7tT7quPJCS2129sDRXzRjpFnUgFbEsd4qy0bHfgqWTI
SR0SqBUS3g3o/gwOw8g8VxE2hM25mfPMD56rBYyHKRpDy3CBc5S/X4uM8ZrBoFXm
fYVg62cD88huH2+ftFddniimFUNMrqclx5Ay23jQc2ABW0RAgofDRrSNakV1HSn3
Kbls2kjI4LRwf6keVMWtA32hVJulofiSKe+NCvcEkPOxVUie2u7ckIJBv1B1kOxf
+K1CpQw4DT3KaXOl/ycDhHmclWKONdXjz4NF4SAnzF3tLhakARyCvmPqcQ9Uw2iN
lu/GnGxkofqxhaKoyVJzku+qwVnEAa7LUdIwRtuC7QMjNmJxdNAZhhN01sjxtUTK
MCt3YcwthzxZXaAnSRESqgFOksTYA6NO7t7b38sLrvY3j/IfrQ0sDNi9xV5v1uzQ
3UXFAly5Dfa1oWqU4tvQTOGCX1iaBD4ctrmtyZeAly1fNKn6LwYCsrg4JfWaW2AC
wH63/xnNOE0NgoVwMQT/A/svluO4CItn5V7qEq+2boXpTJjPWywDMiHSvKb4gPEZ
ofmMr2ru2PZ3ByqDzsVMKyP0SjXj+jmEK3WoBzLeopk3kz2rFqzpoFC82dPlVOiK
ODe5mp9OhMpM+fHKfeMsXVucJs1HuowIDIXiMRWPctr7UJYWTQuTN1xfVfbhRBMW
F7jcSdPGKMW1gSxi3ejcw6pwvcVXKtJgcGE6640qqB1o/5tHEnI47FmGWupE/qkP
1bYfXqsw4bmcxAbjARnseHeDMpNmBMy7/QP9uAmfa3vyoDm2PUqFTOZVWyTp4de9
tA62EAZIm4sJHKOqIp0KhDNu/YXxcNb3gh+hC9wv4rW1HflFwSprDN95BiHY3NYX
0z2v3Nn8JatL0ZFZ88GalGNwuo2Qu7dmkPQB7BmL6OnTGqpJRlxA2dLZ+gqeDDa2
L/egsBi9QJXOLLTg4NDyT3OGweS2Q5ya4plYqfOST6HTRaTdiy4b26onunTdf3/D
sFPHx6bh1X+UvKaQRUpL7ad8KAHPBCWPS9NauyAnSUAOnZAFLLhh2PV+Y0nNHIg8
TiBHnAV1EKgkJR2OuZ1GUtSratBEE7op1kjEl3uAlnRjEdGhXqzqWQGe7TgXBhtQ
5JAKOjzFxOP4POO6a8zw5H8QLo56SJM+E99J4XV3CREfN+Ybuibp1EKPRubRex0X
243Md6fJS9TzncOHGMhVZQuNme1ROlgiStKOUsd3q6YjPB2Q3mWkcqT5gXnWubkB
8ensyw7h1OczDqKEqZOCGPnZUjOSCaLdEPC8cjtbuXDbq4W+knHYDsQlXrfoxTvc
gisww0WBNc9szwkOMDyUQcEEwR7O8PDqE6k+qUjscKI6RDJo4UEMTk1b1EYrPM96
DsMAgb+p5i3LaKOkeph4KPvTpjIWnpwO64PTbc1ebtrGOygNuLWMXJU81hqAopcY
MHKoPYkVKHMmgfK9AWxmabS1TjKYf5UuD9TCBoRygJpz1E4Soi9LTDaj3QSpfQgx
w/uGjMb++c0BtS+dz8ZDSX0RzutmG1VBPZpR9wJ0PTsSTPFPAKeevPG00Mv7m1s2
vnhEQcbkk2AxJQvxf9UD8k7aJ/C0M9oEsJtGgZOLIf2O78giRKqbApyxufFp4o1H
Df1zDOU5UyDvvbWu+4qZwvt75xqFMPvi/c0/zY4baW9oMmfSwZNzOyvCJ9a7daf2
VUtrPJ1oDz6z+yRyrDNUX/HwwSHv0pqDA19Pc7Vi738GMmldouems+1wFMJ8rX9J
TXsYqN/D+r4hC1NgqM8hPf+Arsh4az2+yoKRDxHFwbjqktkNd2gRrBdkioLliRYA
Hoiu59uMt6XnEG8NndmORlZCcrFmo4It7Xkir4kROSBi+uh1BPXLjPTaDKDLXXqw
EX6DSTM+fy3AYj3ovS9lC2ALHLGRGpITQfmxG63VwT+vBAXt9pqnSzfSu6KyS+rc
MHV3cbt28dshPccOnG0SWx9hMyWWYwlCF5Da/mPJQ5N6wu1Rh/2eV8qJbHVdZtQV
Syr9frJX767O6IaOJKJzLIYTRBuJHX6rO8bahlqDpcJWBB9PUQnILxUO7+NGq2NP
r01u99t1h9muFbT3+q+wUfMvl6gOhyc/PL5CoompJLD0+Bfa3igViL9smb5LiwFd
m2P5nIZVDjxC5GzUSuUVU2WVSJ0udgv3Kya30w7e4atR/EPJwVMceagnWflKTrQ3
iTY5BO5BWE5aVdhqrONggrvTJRbrVnp8ym0JbN/2TuL5zlq0Klbzp7L3+1JTFPIS
TYCfwA56y6v03V9fO6FWY0f1QAsWDiaPWvE6yMQLXWJ4S6DIVceauxwPhZbDn2Sz
A/W6HdOjTLUgAka+V7xdAnqv92y9q5WhHyxtgFKDAPq5mmuCMEnG5KZzt5wAiLZ0
N4KRVAyXeFileKqTXLbBaj72Mh42brWtohm2okmM0JuQwvCO6IDrRN2+3lE1MSjE
Uubg2bT1gLlM9XNfJ9On+ijEOdWJpo0n80mGeJe7YdFGAh6taxK0gIxvWva/58Q5
APE5l+hcuLGKS5CuwxnSkOXM6tfZQn9fJNK3BXJFJg914vyInlT3tfNmrAAqzQkc
2Yk7UE5scOMl6T6axAtCtdaY+BDed+FW/i12Lia2Hqv4A77xIUXx4bpd127yeVB8
FK+dMimUTkq0sHSixrxaxlNNjgtvC5qZXhho/uL4LdL4a6zK6/3boIZeG8PAbMQD
RwkY3WFxDrRejJ+0FQwUyKdWEjgByPIE0U3TQw5+VL2Gv/nbMR9t3KipfpfGpK1v
lR+PxGapK86g3BMdQB9uIcFPgOyj1Qh41n+qwVyibmEVwvCdzMWx0tu+kOwRlhLB
yYSPH/+QBN91R7puaNjFx/3YilUAbxKjAkY+5NQd+8BlkGWDt16XF/IAZwzRQa/8
n3lGmVVuXqzgS7Y3LlCNsvNyGn7sYsveN70qxK44kRq0jYMCDBQOxXwRmSxLZU5O
8NjTgCatL8qm2nrgVf0yenO6G1zhLPJKlV5RofF2yeIFfNTadsQk51LpTd+rwrch
yldYVfxkYG5UZQQeFAlB551XPPKoPRXFB6hz9XOMy0GCaJRjqsMreJxurObKWkPX
O5o/vydEKtRMwYnw2FmJC9vuHsuyxuTudJ67/m82Aq3+/QuM0ml/iIPLyJwptkic
XwHbvZtjwS4EUC5PdJD/FJSnonMEfwf1waE98WKIqXV/+I4ygVw+FKAEmVeQfTYs
XAfytRd+672g7m2QnhBN6YcUBiVZ8CjDeHRuIe7lIi5TB9DKDMqweC5IZUvWQrbM
fYBu3tUupdxzTKU2enZp723faD6/NR+aWMbe7LTdlrnCYqlv39HNi/tBUyznGn5A
EQr0VnBzWdKublGKC+FCoSTgf1VnYVtwG50G51MFIRcFmPuOwrYQe/Pa9Pv4LpZJ
gnLKLgQgifx6UWwz6RhZRoEfrJRnS1/b7CQvVoorEct96zZFZVnbmhPqf8QzcX+8
rO8Aa8UJrF4pnOb2TazMa1T4u1rvE/KPN5QlSR5whh0KKfJ70qvryt1o41/6wcA2
qU2ZuIQ5Ue+36M0GqU4iO1TZO9Wz9XUXjWiOksJxXPdV35x3SzKQo+kAucDj/Ytq
fKhC/n3jvWjpAEv5XSKOd2TeuSAfAr1N7vTioOTURJBQkpHWZJdNTES3ctaQF7jN
2No2Axqujzn5tmiedWRZrjHzNY6Vs0lc84E8YLizC+hg8qG/U5XgCmXyYnY/t+y2
oxQIIrVd+OZ5SQowIHsWGf/JY2ZVfxnU0geHwNIih1MRMYgQnaDQ7qf5SdXMiuvH
zxbZAv7O+BLEchqu6jeA9FKFtwaCOSPdEel6KihUYexA1WwgePFi4qL8awFq75oQ
ncFRXNRhaiNiEQllU4PNOilrKg188ROjOfIElqYsNonasFq9bnmh0TdeFQ2BMmoP
aVZnXH/puoRPIQ33od5oBmO+MBDBWtcVn3H7wkA1cis9rjI50SEo2zK3EdIuSzQW
aKtbS4e9qiYtjnJZWzaUR4ixH0IKCOespGQdpH3DbUZbnmkkv9IfbaC1Vu7HCZ2i
KXXF554RWJSaxsV86n3fMJ15UIIXVf4EP4yN73nSxU80vdwEZ1msCH4PiDApjtYK
QUsOPDg3SkO6zG4Rh2mdG2Z12OHXhl50ifXW3ErKGfWvzjdxQPasqzRSPZqieHxZ
PI6wbzF9V0WogxbTv2Pujy+jBqWmroGHyMud9iLfu5YNPNwTgrECj2Ek6z+fQlWr
NGHJzHjLe4PpPByEZUMjMF+lIE3BngXn6zGo0t5rBa+W85qv9IB9eNVkphOcp627
PclgCEY/N9+avk1JxZmpDskmZ3ivBrJX4hl+QwxTBh9x/LIPwlHD80ZgUf+9QA0l
DHkpTv+bemLMnJCUWasTVavz1/vqoabyL3p6UwusFRg/vJ1aByn8j+lGfDUeHjgP
4cV4S8WqZMue012wO9/TDx5et3hcjEbik38VE7AfrSoscfEQb0XfAzo/f8hjpobG
dErWZJjNtEBRomGAVM1n/sE37pQ0KkMuSYHN0M2CcDMURm/c+Yk8aFPcszver9Ol
3wokN3tSQYJxWpyR4KDpkd33mzCSm7KgQFtgr8cia9AqbJeFcyyOj5jaSh/PanGf
IgEMT/2gvy2AyFtT2VLy6CIZJCsT3RQpEL+djQnRCYod4Q74fUCMFNTGfpuG+p1q
HYs5KS9zLn/5CaNm0qWoC+JW7hsxnfm0Kypnfyd0rFw5VhSXzWlQ8OMSN+sgYYHz
1dKLhGkjvwm7BWLlJKN6HVG0Tu2khY8DZbzb34csu+SaQH+wzUnRw8dftD1PsX/1
tmsY30FIO402Oey2Um4r5swkp4niU3gcB3+3hNEH3SZ3ngdY6Bj2GSdAYqiK1sUI
dW9fcrOvouECaMNad/n5Hy+zKrGNkE1/ageSuDP7Q4jnjf1VBY4Xi7AjyBp9lXxO
SL0daherDAUOihYttaAoE2C3sajM0kyClEDQz+XiKl0XHbh5tsqjxoa8to90OFRs
R6XKqBZMXPMZzQmwq1+WoBQ0IcmmOPiCeOQXknlfq6vHucWSlLMk09MXumCNVevC
htsuByucCVQugQ5wLW6iA/LON/hZb4o8UmcRhZvzE1otVYnci34PTUsddANxmB5/
1qQxbM/BfPoTNGUk8Zarqzq0d+l39vgUzboasoZ27nAm02jwksyN5BJjiqK58WWr
vdVP/EWfUFmJOMw09IkY3fgfeBV3b8pImUTwd2HN/38ZldiZLGqofkGfWAs/x6A4
qGmk26kPP0c1ANqZ3MxPGhrsL3IQw0FZea0ZX0Dv/9IlelwTUoGcCThX+SoIWdOf
5fdiGVZjgrb+9NnPPv0Ndd6hnN2sUUJ+Qo2WN13hUo422byQWhCcN2BZTi9uJ4je
b7nZVSFny7S/MjnTrgi/PWHrdFJUx88+aPFYjp9NedOt3xogHCWkgd89+38F4cbJ
Okru0aKom+1bT9K+EZHxG9s1fo3Bh41av5wXE0sh+esvGeyNpqsC+apVNgzSn8MF
yv/I/vV8bpfvBuoddVORRFTYNM+oS0398PLfy9up+25NouEWgAYi9V+Uc6rTqfe9
J38gKS1WPM3Eb1/jZtZMunlcph3iG5KdKTJoAOUOGu1Da+MlWfu2wDQD+VRgsFxO
AXDVzYTNLL+SJouz/L1bl+PCduWVvl47Z2yhloiuoRl5Z50eLcmFIK7Te/GmYeIM
F4cCoL4h4t+qeQsxNzJU1hEHxCJFAhB8+/pdsFnZW9RmE7Kz53J9Vk0OG6yraHm4
rE1eoyQ6RK/zPHTzoH6wQrwQ+lgYP/tBc2n9tAcJud2/m7biiqpo3QmFVi9CX08s
fnWbDaZtLkw7tgDDmT1DMnfBRJ3UO659oVjMINR9d+9fykEt5ImtskJT5jKXY9yi
zFDrh6WHxL/hn/YG0wPmNjp/yH9VS+kEkjfWO76tM0tycou0J7C1eTMiGOpY4kM5
suk696Ro+xHGgAmla4R7F2BE7hS1opBUSrq2ZJCQX8IbMYXkxau/iQaa8q3L6C3o
N337cdfXN+5LLYGuMtm269EmEBL4tQCxloVTCUDmz+gDiLIn8mi7fWp0WvGxtY2E
YUidff662FybtkdSo6+UjSQZuPVbpg7bNdUrZziZDUTWWzSfv2zPcljB7xfczIj2
eCS4hDeyFgSeTAL2Pru7JU0u0enTV8/Q6heHxnWp5TQ05AIFLEe4johTIRetb7ec
H9GNRNNQcad/Q2oLS/z8xA0ieLmaTDA1ZiKJbY/WbALvdchmeENhfAIAwf+4p+10
cJyfiBxXQNwrUJOBJc19q8JT3CjknN54fe/9zStlOCvuMLIurdpPvcEz/ZYY2m0b
AQ1CZow0+RbDQPQsF2lgmb+amFhinkDipIgF6n6Y9+dZauPLxDpiEJf5BY/8sEV0
6cWSrtxBGrnAGFpqOrkoKNDtcJ/tduJLi3HWLWmAyN6geTujBaHWCsqqYtN+QjqY
Q9DCje4BbnsC0RiS9PqpAnuj3hbfQWcKvCAgQv6P7CyPjl17pxGq0WWPGhZqCTUI
fmoSwLMm74RHGSVW3BXW+UT0wmwc+OY8HzN45pDOjmAEbeTZdj22wMENSolXa1Er
Ny/a3OeHPbUnCF+UhSYBT2FzdlYu+75fb2qNzY/r3w9VFVC3b8Mr3AohtMVCSAj5
Ie/t3MQpKzSaPs1TfS5yRNKgOzhgIJbSAwCJuTPsZWzaSNCYdQlHKkzb8Wr4IfqO
wdzTYnQJoQYysHZ8zhXBQ4U8EkAVkP3PcqSnyvCsiMYtvf+jOTxRLcuKloSPtn95
4VwsuUnMlEIi/9/V3ll3nAtbcDzg+L8KJ6BE1V5LjMcRT9hgnRruoOzqW9T/n5U0
+eprHR3+nULRhreGMLJ4jM1q5a7ukO0Er1ZP6ij8LyjZgtJqd3LGtH/3mwIqv2IM
rSHOiN5qjTJBbSs+5jmkI3QLn0HHCfhtYWhoZKjjc+V78diz+jWgvorNJ0TZXRZ9
gq2ICYKAAKEBl2qAVOlUeDN6Hvnw63GodUyxS8Yb3idctjgNTkkn//NvvxBZ9kAQ
TlR5NP60JTYhtJonyJd2pzw66xgQx03PfUOymxdxLAi2N/6OCP8/DHrdc6MiAPTF
WWdPSdKwGLIu7XY/J/no7WCJFyQ4l1FGxtO+1a1LV+2keueQyqgnXxXP6dDjMR4D
c0K8SNocnEIWEPZoQkW9u+eY8S2zmCqEhCZZDDocrqZWyMOyMD1syOPy1likhh30
zW8Qgc+6e+fDtsoshpRlWCJlRXhWo3Nb/VzxYZRDf7jCfSVMPOdxWTvukS8swjiW
oTGZb/Sj6w2oXCHJl3L0ytEoMvRUMLC7KIH+TFcQRMgnWGNpAANZ8HcOVhQL9AEc
fu67L2DfKpENqGymwtz35NUIM6v78xFtP6sRL1KmdB2RzPJqDN7VRnKFX7YdBTkV
obEN/Zk9VvsJoPvhKmZfoHTqWytTknThUYFG3XY1S2WKEUGWYWUuZgfXC19QHNYs
v6+4+tvxbKD28vuAbKC67i+O43Tp+UA02Ps1mZefkbFHbxJHPNXFHibWSC2T/LWG
Rj+2e4QLFy+OUIAZq6EfPxHnN7fbP9HHU8eMVahiNUurJgEVbjZBoCYZMUEI/Ob5
sSjhxCHKDg/W0Cmam4vZnVxf5sF7pQ6ws2H7gLXq7Tvi4Oiif/j9dttJXgI9HDC6
gR9jk1D/3yntnAa7SbGLKFiEpyJRfjzO94DQDlDF2Ixkh1bSXNgL5YPnQ6PvDzvd
UIKaZEeTkzDkG26fIBqfpI/ArBAAKTsV4KI95fNjAwJideEeDqPqW27EQa76aJOi
bpvTAaF9DOn3pB+yjFKyJsMWDA5GyZClsMB08Y19JRi28EUK6k1/HWTHHSQhL4PY
J0AMG2azwRChXBHucafPC6nxPUQkVvzbhqSIA6kfYlenk63d/k4/KAgCPfT9fy3T
FHC2BomkIUyKfh6DGkDbABqqVnfWKId4g1GCKDwsqgXdilYI0nk2r7Ciee+B46Ty
Ot/aI7Xl3cTTs0w6n5ELrlxHc+UttrgDefioQZSMm2egJuNMJLwV91ONezKl6bkp
9sfozezMb/0s0N3z7Y17/BPSU1Mi0ZmUdO6b8NZ3cojHduk9mH+bUDPKiNaxO1yS
qb6LxXCuTqdnl2A99P4bGRtTA6wWB1T8+B8Dqe+bLhTN6TIYzl8FJIWDU1VJHE0f
cA//5E2jogNAdajl8OVm97DmxYY0ADfVYJYHpaSxwBt8WPDJhvpgQ1CS/rAlT0C3
byOMpK55KOcYU0tn+Vo/zc49x67GwFp8q2SInaiTtIDl8dgSLUKqepFK9UBxZlV5
YfdstusomXhc4Fot5XXQLi4lXPG13MZ7+37ahPV815p/IQuFKiwm131vJs+XhGBn
zB/Ak6yZvqYch5uewoJcQO3lG3rOJB0hKzKFN+G3f6l5PYgqNWyiQdATL6sppEn/
YlC39Dr5mPTl03llt2iGkI3L6Z/mZEBRQizC74RHOqHqoz/fx7//kV2m1wMomm8S
6KCeBil6+r67TG/aGpLjJGaT302cI/8XLE/PGxu40aJJDOmFVhcOsHeY0rZwAHI5
CI82Zvd7HzlmuGdw6uyUO9ykoztiTadwPOed73LLF3DTYWVS78uEqrtkqX0iFKF+
7jYKypPtKtKfHjPHh9S9bA3aYFHTjFgi6CG3mDhF/3b5l8KY4og/pzqXhbgIjJ7b
uDZaGMaUlB9YUo1s6OwjLxVY+MCTCvwJJHjTljb7lUu/ha1vzXanegev44Nw2yyy
+qJfbWmSrLbHDi99AIW/Xbh1ybzXF2kdQYPFcW54zYFTRWsHj8Reyu7wYaR5MfKo
kUnZSBEorUeSFO5LqH/3n7nUV6UMcFABYohn5w4X/H0z3Cd0O4/yfNFzFrUl0eV/
VspYlENK5z5DLrBOMTY08sYPd6lPoyr443twn1w9RJWQMlHYZ/wMaQ+5YUO7wRe+
Szyvvd1GAnAAexPZEcMx7HAoJ0zmcIf90NCHbUkr1qo7ladMgpUa+RHIMDYOkZwD
sy/EBkWetKhm+9xCz3TFAJuWXPD8y4/qh/xn176BB1nxERtOCo8SC/siFlCvF+rC
j7gtZVwguOBxeflO5E6+zFG74rsKQnb5Xl8lkryzVXwZUOqzlmriyGeofItS4w4N
8EU+xa92OGFuZ4OaY9AshE0UVjyKpXt8xbEhwpTnQUplteoZ1XIsK1mojJuOM3U1
nowpUtHRbKRJ3ipV3YT4LYDdC1VDM7ce0Ylg9vvNy18EAYvHeL/qR6b0AJ/z1b5A
CW4m3eVgkGRk/dd8d/dIZloUN1Sj/Qwd7fKVJkItR7o5R0g8iFP19rbJJI4XQvvg
8M7C8IWMsSAeesRAF/bnrik+Nyg2oOcNFy7lpCbg6m5ycmwku3bf2bMcf2NQVM01
wQjJVJZDJw2YlSyNRe5Smh0KQ/ruocI6kDOHHOEnMJPDMr+dhS6A8+MwZZrcVZDD
m3O9IVZ1iuz09nFuoagdTJMlCZ0nJCFdel1lNL/edz0MGH1sZkJA+cigjgeUteUW
zzgfFQv62KQfn1kQKviw8xvS1HeVc4Z7ZnIy3BeFzZqoG88ie6goRoK2WP50W3Fq
HTLJd6orObxyRnw64hDKzNbq1tKPW2nnkXgutoeHv295d+BYuts9YRrA0jrHSq0s
7v1HoZmzRGB1s7pXkIFTe0htEGYOEyTdYWOH6NgyCsVojoZOSILMFY2cQ//CcJGX
op8HtgvK6bk3ueLUz2uUt6KvV2BYKyUazVWmIXEbWe8RVkRsW+Wghw8iwr36b/ov
/wJtQz4cngRtxV5VU/wzp0hzaOLc9k1HZrB6sMxQ6broRfIFaInZ0yyRIdeg82o7
aHOuguWDw0Az9SU3m0XkZRS9nhgfCCFQuD1ZbwWUPcI57376Xa7xnU5Hl/40iGEs
i53zTCOCzbMvULCtEiKhV5ADAe/fhCgXqRNnpLKN866Q8QK16HkR2qQO5ZPQb8ok
wCtjaftNfxx2/RVL9bX83FElvU/Me9ck+mqCYPdaVtHRUE0P1vBwC+G97yWQ9Ejy
OsWE5SIhDM6U8zO9sC2m/g3UBzOdg5+tzc8qojFoZBkiU+6NnNGx2n1F5/F27BWQ
NWPQaJ8vrPcTBUQJonn9mF8A3iRYJ5/pQDlgJTSXAe8jMUpFdtc2/pIGTQMQgamT
qLXhAlrDqi0clm2+RNFpzDWfsnXBXsS02YBJRfQY51PPn+TPbf7NBEGLX3lY/Yqy
spG+QQ2ty0I5ijfY0Sm1k2UeRL1k0l28HusunAlO2owZOam9w+KGwtcbcPUX82p7
f0q6iBlt3GSg+/2wziP+PGCf7B7Qk+jXgJBDba9orRx1OprsdSUeBn3skQdfcTUH
oc1YSxQ54zYthMaGvZ8606jZkyFgrm9dU0xv0oNztKCTX2PvPz6xbzY0wN+dr66Z
22ybsvgkL8BnHHeviySM9rHFJ29AyZ3A/pziuat2lk74YDTSY6oAUY+Q2W5gnhvU
vLq5hcvn+rZZ4atsLuUgJ4sUgCfeYXaguXrHItAbASqsS54l6ui/xfTPMbkOCSgJ
Fz8nLEWTNgwxJKgP/JT1cT28JbmEoLGoBgP3ov/EBUSWiRC9Rfw9kSHZ9HmGbKnd
YE1u5KKt0dNQczPZqYv06Aumz1J6BtKctq9uEUt0DqTTNGcC1L7khKPGKp4p7nA3
7oAt7cYky0J1Y0jhGc3ZVQLFWIpVdh06zaCKU3avRxTY1a9iGTfB0OZ/1L0HJhta
kkbTVerIBmmG0OmoQyUcaSijWJAwrIsBm7ruCSaLWCfyTsIebGJ9SHJ3ualyImdp
qTmWq00H0d/rKiWKf7Yo5jquo5kcULEQbaWk7y2tfkQSa0pDm7prWKphDEcQpyef
tRdrlASNHap2zXNKKDqqqkvZ1CJsPadjmUWLSxsO1Z/2GJ5f45nAuc00YMsrqVZy
vWD0gyS+d8uWzBzTYf6W33NSb178+WsL/XQ/3f1g6StLiBKq5bOR81YTO1u3ahn5
e9+DadDmyo2d7jw50eyPdeGZttsgfNq6HEjNvY/SHfBymYBAvxJdWl/IrUgvMxXG
QayiQcV3HC5n8guenVw/n97Xyl10HUT//IP989qE/DAYP2h8HJm7bSQTG7D7smVw
Tqt3KVD546XzlqC9uWSRpiySSaZHdac2Q/SnYsg4NOqsa8BxXvP3z21p//ky9OD2
kU8hvLA50ouIG/qHELBWgZ8sPLnHfAd2BRy+cuqZnVHvtZeYAh5cJSDGAfCX8p4I
2iwFj4uoGaICTf8SknDg7nBOV61pd8fmvsv1WBUzenZUPgnCeiIjfyhw7apqODeX
aVKc2wzKdLnz7+vUASeGdmFFw4gu8gb2CpVfpNNWRticaqwc5yNqWSZoNEORFpV9
YRN5/jSgy1jIvm3SPbL3XeU7Lccbipw8OPtoPBP/nT8spjb8NJ3ajNP2Zt5TtSFs
PvBhogakzAk6MGTtL4Aww6JG33NYd055JBUyzY/2sTQGjbbLaqM1lo1cRZelm528
o1jDEqzqMpXK2EZSaIZ4kPrRz6MvYDzIq+1rDcDyCSL/8cMm5WdyYsyR9AwpG7fR
5ouEzpCSHZZKAzIVygUuM03TkYW+wX0mX9NUfFyDvpAkNTibBqt5adkCU9AE4Y5E
hT+947u8F5mMULc4cTSjA684VzvoMi2Dj3gupJ+PhBhb8jwmxMHLNKSUJUcM0dkl
WOtfsgkLZlGDmLV2JQdwdjFl9BrcuzjcfOpXQm5O0TTzmY2s1mlHX79fUXwWCB4A
ccwuhANMuL8rEPMkgY2e/JvrtWZANqilx2TJAWqVRz8s6/YLTU3eB+ZgRcIaBbgd
h2Kk3iE5VeREVChYCL5urLWCuyUODGAWXw38xEIbOtmedkKGZn2R89NFH+Iv4Tg/
0I3w0O7sgVNL9B3qwtpdhl2BGGnA6T8LmxjoWSsClBC4haJQINt4Ywy9U+UB752U
SBYdbiqCJIHchTat4hA5rSRl59KfKvF4plyfdRbgxizEykglHmQ8+vc/vGowIm1/
2vbobdcRXeecJnSfMQKwwke/5u94U5yN2cXA5oR++LGqPl9DpcumXfUw7Fl4pzRc
/GFDs/5Hv6bcu2hUbk80BAAUqHsDm7DxMbW79aZ9mrzaSdXGY9hN3qBOQRSM5CpY
SsbFCfV6A9Mw4kQRdLlVw8bpm2FV0lrfp8YU6/RfG7N14S3zSNOGPXAsb0L3+20+
+6CksIEK7X3l+2LhzOgsxCBPpHQvhqbCvwM1JHfrQypu8/Mn0K5YUeUjmVFSR9NX
/BpWNJ218hQnspqHBdekfsBAI9jAY3/hPVtGzuHjROzrph19RoBpuTHvrpVnWHP1
NPgkLj01buM/vniPjBF3o2t9v2bWFfCfEFzEjJI1GGJoeh0SR3KbZg7Bqaw8XT2Z
R82YYHTuGur2xsQUIJZn8nXYMJNgQiT+UqY8fxS4Q6jAmUCFDbZW0FcmKJkO9EBg
mICNCrCWCBhyi4f14sBkSBI7y0ztzmM8gJq6gHsrU4zk/90+n1MFZIEEqi54qovn
0w68FeLkrV0NKp+SAd6Tn3gBgR1GmGBu+tL5vpH97k+Hfe9LYsgp+XQ94lbKHbeY
byrKzfnK6ckiJ3D6AEWwaqnNP85MJvWnKVsPG5RRN4bYJQZhZSmmbz8ok/zszhMz
ek97XrMGaEpG20Q0AFx6GBe9uatYLBgIjyzIAHN0cxI4zbPt3ixWzt3jVPZlSfoQ
wJZ1GtP06Wwb8EUG0/b8J3jkmf2sxxcrRQa6O8LNaW5roMQDIuLY8gu/Q1zc7kLD
n2chNOSSWgKuVhvWgN/bEC+UPoOS5snICmMWo0GPAETohNGIafbCD83hAtiFieSF
283ebVVu3YLVW4tlpCThOtWinHwMqnrLhqDY26QT29MsW8T/1x7C+SVytnbj3UkZ
PwxG7Ym0+35qLTTCdFYjWTvuI4MA1xK7AVk+1GUFgtaa+Y3WR0BOpBvvPZNa470V
3DVz+hy9Df4cxIx8tZYGeE8uEclkojt0WVM1XmxndNfwrTnwdpWxC+/8nlW+z6tW
thl/3702eqekAnaA77PHIce3uMWpquMFfMQkzih0HYsiq7TBVyeWriQoN8vI18bO
rkvk4Uyd/XfD0xBWtk+XwqTlvuhO1mvNpz5+zO9EG2lIb7PfekB4wg/YnJJPjY82
xgBxu0r6EtUIuIF7fQlp47qtbhNsbQYJ0QAOp9CDf4ngLlMUp9Uo+VjQN/oBXPPf
Mp5ZYtcAWYWHU5UsSDNCmZh8cpUVSTA1QbOmMDWMXT6COvc2JMunapgAoZK3mEMu
IlB8v/yXvvJ6KaCMUlErsPhc5P2+189iA9EHiOm+nIc/Oq2WDibctorCBh1pJPPn
bfLarZGcoRI9fJ6lsNo9uALksuMuBPXCBLyEQj+A4W5y3w7G7oP/tUW49/5rAdxl
kn87n2utOlVyLl4c3xcpY+GYcURN3Ebh6fK/DvxeMrDAp/J4q0vg7MDZsRBpNkve
4jgFlPlPN5XdKiNtVH7vSOkS0JFNGmwX8z8jM9JR7Tefb7tnzSjZDVBAsYNC/hfK
w9eIq0461BPyuy3n4AitwiMBlKv70WQKFAz/hPLWOyovN1do/xISswjjD7zlNA+6
g/2T+KEB5aPK5m+gKIDMcvozTOO8oBkGEHYbqm6PS6j+oSm5IqLpxaQw2GXfDdTO
cEo1tix69rRUDslPupmDFX7CS1SsZrDIFtcqX89nhH1qD9WRkMGVc35c2/0Mt2em
J9jDUv3UK1O6i9PpAAz/X3qH5VmLGg1poo0S3SFRyK9DXZAJr64SGy7TXqv3BbZ5
uF9XF425EgjrRqzUO5DIkHRqWXk6aMQy0AbdDTkhTqNuBi6jo/xrpXSetogjapFS
Cq9N85X9s0OP8iJa0aTqOiArTCVOrPS+JkUFe5UG5xG4tkecFpPcEEjSe5pNgQoG
JM4YtqwgXkFdrCMbSE79Rr/H8y6YSlOnwQh5phdmH3ZyescBDGiBkL4QCMQSmr3T
c9yag5QWHtK0XB1l+vqUea5THug1DnTlk0+yDQ1DpVGmASKl2GCuKpnJGs4nCz5s
HP7MV9TPfCrL2/L2BbuC9MHDjYo875ibN0MIS2Huq5SXwLQLgEqQo6ibNF1icJMB
OO/LuIBqmchOVL2X4mPOmdHAqio9YjHN2jEy18hfUkE3DsDSUB50tPbmv0ypUN5m
nZ/c4useP7hSdp4dJKUj34gnthg9ezByDxA4qF51PMuNA9xlEEImIa1b9GbY2Rql
lOkGLOaLZTtenq1+7M/TJomnjo3KTaOiXhrz0d1FcvkrE+xQbDm7p+0+1AlnKoBn
5XFXtStYuoDxWk9tNzFW9I6nxr3cTutsBsxFw2mrAfH8Emg7E84KFCiiR+OWRJep
RI1Y73iITEhjtexbwmmqqSPCrS7QoYbhb/2DX5Sid6bNxYLqcHywXpe1xwCVHlUa
mo91IeIRqY3eJz6WSqOq+Jq5Juxhh7PgUuh6F1a8FERyOwYaO3+x99d9uiNmcsHT
3ozqhDx+Inpd2GMRk2SmJnZdbligEIdlIlGGXGAgw3CikJSQrMFEvk0Ab9rQhpan
iCRpZ3Hb6V0nw4i2QhI5UYRM4Gc8GPLFzy6WBiP1k93j8Jp7VXBPefABnLTqQAzn
z4f7vvUaqMI9ky/jhLGCuu1BwU7CSc1kjAc3YobOeV+IeZeW3sr92CoFX0gVcvnV
G9xBpBDjBTKPT3PDLYPUL+cpkyGz93O2OZLMfQqOUrMlHfYon5sgAv/GuUxo1qj0
A+1ox0NH3z9k35fun9afY7OEvoo8ujcjtWMyevNDarB4C00Jj1ZRohqi4Zvfav+I
s6mlt5oYxTgv7BZncQ6z28yNx06zifNkWeWNZ3nAb74bJK7a8wGAcPtO0EvGuWNO
n7fPBv6C3x1PXKRLSqe9XdFsyIYkDCZokgRQ/WU+iZBv59oQkjJEs+JdzzaPodzT
PiFNgz1fIr9HFU2zJCN4VqSio26abGUeLc6FIMKnrbkp/FuNmC8kfGjfDx6v8qkf
cIxQCk17OqCZasrvjy0KxIu/rVFYhfZrHoT5guk04R4K1MtOcReLiuo+OeAHW2jY
tELGNJVjLtaR2TbDxXsyfRdWqnyfrMakWu45KRtbrYG6EGNzTTPAVAbxYqbH3q4v
MDyxvov+UsxJKvRnvAZb8hvIsqobYvdzbrELz8TTCu2jHnFE4jhNKo0cndQNNXR4
F3CLdrm5K5tLmLoBjJSWEVnsHFtcg5hJ6yjuLhdIBgctSxGJhFWdRKsZ5RAwB8aV
U9w9rrXkNhmUcmCz3mv7KTknPV/bBeFZt/AkqCeBG+xeRqf9ttd3trer6TOpAt94
S6Ey7Hy8VOGDP3UatZ6qbpLNCqAgGTu0kDGLiPdNZCp9Qb8njov53uRNj+t8y8xM
7Xw0QHoFPmdBTtdUlVqoVIHFqG56rcIx0SN3NEfKFvf3CAsrVNoAJpUzThXq4X3H
WK/gnv5z2Qo//BXWOj8WuVmjZ9w6BAnYY7Iqa+rcqcPOqEkkczfYMPSwIQvfevTT
oloIz3H6Mk3xNvm8tE9QIso8OPAlHZEtxpDhapcHrJlZAkTwhNuTRkungmN9c+FQ
UCN8hOQk4e40ESog9NGw7/XEsVBVue9lbCFA3SeA8vTyb7Ze+uD6081vCHRkqoKY
7Q3G3NUUPKFHZzfO0HLdtiokHX4jKtx8msCFTrdV3AIoxEtuJWZmX8eWfZdAPh50
w/M6TtcPTxOxCMxmDMA6Rga9n6vvb8Lbzgc08piAO7cQmisyOp54jBgI7BSLB6zg
YZcfNT4T/zJ9by4D+0GdN8eaPnfAcbc34iuSaBjtPW2R14PBp5P1KkU9xrKvmeex
vTUMj/1UMgY/oe3PZlD075gA8f3IOaylJFcN/FfhQfr8407K9hihcOyT/bUdjwrb
vxEE6WJ8neE0vTsaMp3QJCXtSjfhYMzbVkcSNKvaC03j3wud7sL76M8YEP9jpwug
fMeJIw+sJFJSTaeWFROiAREogIUejjZTQBmSI1G7A4zZCh37ls3BR4emFFO42MtY
padjqSHVCL2oMGl16YA//TF8qvqb3JrwaP0LAMNuIh3yvhITEdll0W4Cx55kSpIO
8QuN8AwgLSXzb/BlogZfDYTSopsGlXEBjQISsEQFzJPmGK158VadeJTN6T9Kk19F
OvpazU/GRVLCmSVhc+aWyhgonqL65AmKK6w86K9YuhkzeF5PZCSiTMGTsa5+SWpr
Toc5wvO2tp6AnYpex/+p8fDHCRwoPT1VjdjDW0WQK83lMrqNsMCerV6RDpklkQCd
au8gs0DwzGNrAcFsHlnKfZsVGnFiEA6m5eMk7BdXj8m5ROuCNKp8wBZElrxGbZma
5i5nExDdaR8LuOTxvs4ou+HvsgY0EmbrrU0yTcohsLxTcMS545xxs9i2SU8PU93i
Azci7LQtzxjiW2GeIJLm13bee/xCp3yH3d0/yjd9ylFRgc2vejpfKJOWGioviPTG
6LhlERh7OLelqKHJIOjWYnUQFWEGi86aA04HN1Iu/CcMbkyZfGNkBuYFGWHWS9pE
9NuSQgTLCi7sQfw/1mEehuvHGUJxPMacfRve4f34oyUcoflLHlaeSFVWSfyMV9L6
bvqoyjhbqZXjDVcQjphEBEi9Pro/RSzj0JTtQLOWZBi+dGHdGdaRWwqOa7IKlIZp
u+mkERHVs8AlMMmD9PpvE2eKatmeBJp1z+echE+lFyu1XalyzYW7KLhhxgrRsytV
eUM0rh/23wtLNZcxqUK1jYIDVXPhcJl5WLsX8lIML90LUeBpipyHHPxY960Fhk8p
PNswBO6tscGP+hBhvtZh/vvVB2JgkavBq+G4/X3H8OIAqViCH4uU2OpFRviX1etL
8QyTWIsmv+C0rv68RGmE8PPUDXUi2fp95h7oo4qeUdqbkMwN5DELyhVZHUEQwA6l
3mjzGcI95d+GC1xy6kVj4W/ZF+WaJH5yi/dlhLoDjX4tS0ikUvLU9dM2VmuAdlAQ
cr3D9TENWKxVhiAmi1q4Yi4JGHhLEmH3KEpFmHDNPIBTlf8m4YYoZdjUwxNMMTPy
817mVH1jIRHt8tXI5M64uYgwgzI1Yxt/7pfXrANhVpP3wz5UbZnUiMbwHaFegcsE
8ZppW0KteRXlaCWXoSa5lA/Ig9FwZy1jWNLitf7dF1rM1cXosq6gLPSyap0tw4i/
eKXMXg9qv2GjoJWvF0V7hFV5kX5hFhP4dIcI6sg7Jtc8bS0azV47y2SHQD2zyo9V
Rd75yveQhOfHkGI2tIKD4O2984LZuDaC9yigMnBOLs+a1VOmdhCmEA1WwLwfpq7E
fKoVFxFbijbT2OG3YHT65MEOuid+z7qRlZQBdiZiFd6lD4dm3igfQFrXFIE2rXCd
fIloiErpWMuOr9d90rcJM1N9YoKUwcubPTq6rjkrNnSeAXFKr/D7tVYmka1xGSOT
MJpkup4aTFvTNCRUwJNLiC426u6q6q+iWqzHCkxOcJGYe61QtbfQPXx+85/MMkmd
kGzlCnE24lRXCXjDMNgjqkB22ufy9YxOGstfIHIaROkOtssWrLQvqkD2Y25jLjjG
QVXfQZuvijrOhp6DuRFeJTDLFqnfU70UqeYRgNqsrUJMSlH5bOnSwW1UnmbT43QK
KNgwMbvnKPx30yD2ySpWG7n5gPPZ1SpRE9Vz+WgW9aqFNS5ifGrvpXaAynL4xDTN
7LJwOewTpDZWNtJ6MLkRm3kbW6WV8ZBmW81Low5r2E/QrgsVnPSaftNfZDedPcSL
gXENQfYDJDWbuNYEG0PtsnmOrBgOyIKg3kmtvcMhtXlCd8Rb+WSPmNmYavydubPy
6hG1lB1Cvj7mhJrNROr4nkIG0mV8Kf+eiilXggjgXyHLPQHJptB9dXcRuukyjH37
rVXN+qiRS1vb6MJcP65Q9VVuJIiepgdoM1ZwQOitGRN+eI5q4/ChzJGD8BlFhS3+
KFATFsedmy3PvqE+4hli0kjyp84SXEU4TSleBFYykXvMhk+w4Q9ujhfngYNJJpM1
XQM66KwYNNZdocCLUx640ikjjU3bAky2j1FR51/aRmUyWfkD0BNAwXiMZXzT7bGB
D8dCdTXstZtTRZ4MYM2aZOlTe0Lu3jp0okj9pT1hEVx6NIu0yJ3arrlleK8GEiiz
bC7j97r5FIyhpewhi4zlngiFUH1Y8EjqaLeHJI5gR25z3mxF6twOETEjTs5HKaHE
ZoBCp9MoEn5Oz1HTsn83YHdxXUtlwznd0qNR+k2ITNlUTivJZ1A+v4JZhrnlheEx
odwI7ggpJs0wYiMkFuigBV58WD9ycTFjjM9HeOXCRBNwZrQiazJRlH1vaAINB9Z8
7eKxv2j6BGLFPIiDGkQ8BJt7yosjMbQWbT6ZiKtmRn4Jo0CPrxPte0XRjXGgbiln
ickMo8NiCV3ej76cakbNB62vCmHAeWEoSJAdyppCVaPW6mI1LxN7RJav0bRY+0EM
l0knAzL0c7zLQPEaB5hrJdZUOwz8E7QoZSFxdPeE5jN1Kdx0WCau15qZn7V93c/D
uuWDdJq7RD4CtnWVFgGmcsUJrzzRUROPZAnbuDkJPD9YstXdwu9qnTBDDjI6On00
yObNeHmEAELLIV/t0bJwcc9kdvI4OLV3rstZkJUvw/9P3tBxYZP+G3qJUeFJPTrV
dc0BKcmtciWfDK5CZFnb/BjTditzR1QLo3xBF9/CWU5PSbuJDZvHRdkIXgDIurjg
afmsXDpsz42lIdlL3OztNZIfh3m0+MzmEHGB5lQTUU6mdC3+iG0AS0gUmB7iWYPQ
au0wKhq+gQUFQP0qU91SKc4fH3wx4Na7Lqj4WIHe26GsNkO2TiHLWcx4CvqxzOvG
kMJNAeaghGqpRHh1g4YzHjrxDDihcQTT0dtfb4gt6HhxGf4XJchvZ9sxhG9RMV0M
uogg7rDxbt0Wx7dFjq3R0oRndZ+DGvOyfzOkVlpdatfvOdwkIc8IMT1Hsbe+AXll
pVF7MjfDtEb4GLVPHE3QOtEP9MOcB/lKi0AqF8Tv7vhXqmMJBki247QaA4gKp2ny
j1s0mWlGVrWbca1DtlWCJ/XMjT1IYPkEzLkq7MTHargs5oqXM3VRlIRlKNt+BS94
e8bnbrzAQW8qBoYjDORcnGhkX0UzpjFIM5SD/jGYNQrOKJn3V6fusHQg09lgpV8B
qB7mToYWXQliSYqi+WVdql94zs+ldOqceGJnHdIZhrlcrRRKYpebC7xjEVHNJFpy
ycC4GlO+VpttNLLJ0/9Aw4y6ZIeytW1v6AtzKGOuu7XeE6aiWDLAbQ/XaUToH2Xl
XdnX8A3b8Nm6pwlN1OLxQugXh9xApg9bunnEbWqaX2MD6SBfS1bGdS+XN9slrmER
0rNeUEl9fB3mbm1JvDSLwD1zzrPl47elm80aNgEq+SFraDsRX02pOTf6QH2YQje0
8Rm/davzkzDHmc8pmy7rPins0/y+WyfOvz+58V2yy34vhxy+NPOE8l81Eg6HJuc8
W9ZpudZ2pcJ18XPJqWVJTidKgxi/4220DAomz0QxI7Qp/cgLqEPRd07YFx4TDDWw
B1xfaWykPnAdDOfDENeo8BR5SqkNjj04mwkG18OaKcZvRsCOR1F2uwjoY1nG1Lx9
z5CJW8kI5UamkZTXckv/JaZop4ZAo1hgcbKYqOt+Dt+iRNI+QLqV8a68RF7M+TFc
bp21THj4P/5QockTTsWXEZNCemV9OMHEpq/D9lg5xtYlnOZBz8ZsXUQI65a6c3Sl
zwCcJn8i6pvnV+W1BX+vqVMeCtcamQ8E4W7gxiWDz9e6hLw7lEBOTZPzjOb/Ju53
au0w2QKvBQHXmbNzU7JS4qTcBb7cR4rhUUsfMPv4Hs3cKvY0AFj0MhfY663SoI41
e9N/w7aD/bKb9kRKJZHhPkPrH+L0iHTU4RlpNKDnU6e8hc6X5bZwImzucCKrglKu
AhGfPULWU5zecLnw7HCNn4dFoMZEXuXk8boGurQ8Y48BhmlIa4l3PmS6LxjnfxaT
IHA7ll+u94dsKvIsPb6fF4GYRtn5iCa+zNLzTzJkhQuWOkkl6aCRy/SlVLIVgp/V
ybkjSfXCiwUC0JVnQu+xsPNVsV1575OmFlg2fgWEQY0We/U5t3ztV/OnB7Fyo1AA
p27Pm03xBXovw3hqZRGQoSFW/xFS4YMFp3C5fpXx746+0xs3v/GYyt50w8D95mjU
jE6Dyt7Nv7+Ue4PxPET8lKkrekCzf5UzFyPwcjkOh7XsiUmAHqcFbAsordgRlhS7
k4G12qB1aBN5ZwOIyqITLKqK2t82Mz2xoYNaQ2Yj2VQEBKH04ggzD49bVgo4inlN
s4KrVcoj3Utl2MNLUuOwBaUmxQETAktxhWcNsw1rWhjBdPFaU0ww/sKO/eppfPX7
SRxz38lrL0tp6cXWH8bRaI8tpi6dYariHuZJnnf1POLZGKC3TRNu5514mZK+dMYX
3wRNcRMjU1K5WK+mj6bdBLQK7r+hEZ8tWqPPaeQEe25J6AWZ8EbZaVhd6pFGb8eB
nU2svkkomIcvHWKwgUAzgsyx+XdYcC2eQ05FLmCiDnC6ccENeehc8QaaNIEYZGUr
haCfaWtbJRnKd6q+wMLtxs8XeeYi6qa6JYd4ZZrr8x5bjP0f+GA6YgF7xYdQ0/Fn
Q03kJr8egW9W1SrK0+JdV0TA0knnVq03N2QAFL3JvFWFpOy/yBcaBIep0qrex7mA
5nAFYtSkYIwGvgf+jbjc7k35Q3cLYcVkuY5sO6qyk8oJBMGa/KPJVS3kjEq/V66z
JlifTUfUj6zhNjp7pIZAf86+RAtL03hJjelXI0yS3SWVT7s+brxe1umMd2Vpgk+8
kAjvslBaWdsnxlEZRLVjNIiIkgWmdwQbnRpGqFF6sVHDzz+tQoa0hSZ95qFX3ICX
B0zvcWD8ckGzrcG3wNTuBla6h5kTlNeZ0VYMhMlAnxExjxoWWz6O0cap3r9IkzTg
TYmqz/583HIKp8T43ezXTHtc+RQCa2kVbWMj+8urmI+yMdGfHPvfr28oiFH3L1YP
eoXLgihKSDBGBdLIhoRc7ueqyNkD+D3UlecwhNJchZEJ3yz0n4VaW6UgGj/l1gc6
YeNAYgLXUWYY1Gx8052iQxoYy/XMz4QDnUuWi8fHso4PXQua1Fi//nq1uJiOpVWC
3A/g5QNRLlmY+hBtgFMMMloOcQnkFLOhQINLQ+Af136Odiv576mQpa5P6ewv+03w
DkXLiaysc+VWo7SPTkdMx3AyYro1Zeax0lg3ZP36VqQJJFYp+8FR30tvK9jIC9X8
YoEjZXLClLWu5J6ajhLAt7toJd3oaUPsInHcO3am4E6Aof3xVXjtBMemhDeExIqD
40ijOSqupccE09eg9WeMrcnmtOCYU3q6uvoFsXkVlPyMlVm23JQAsZdYIdhPubQ3
t3R9QPC5p41Hp32OF5qu5Xhe22aw6GKVYZ+oPVPh3TAasMO53Z4hQKHlhXm8x1ZB
XG1bqAynu1iTlJVXdhlIT9AvFAmHqcbtB9i2HPKORuiP4PnzFuE053xe3OP+sG7G
mhN3MVDz0Ojo0Pcrl8uaEDgge6/dZT0ecuS1RigoIsOlF+iKjPefBSf2r725wEy+
WcA8aI04KGsDQImOGoRBsZ7P4LM5cN63mXhgImvP64yaAS7lcmBqbPdgniibfWnI
S2xeAUg0qts1GOuWr8R00GTdHjm5IYXd8s1UDALEYCJ13sJ7MCRaw6QBasX0DU9S
YfQD1HMTdJK2PIV0FfnDkhGhGAbFwvXqD3vXSyLD+7M0bID8XiYaWbOei15WAN/O
bsKvHdW6932O3jZpajvfnQUIdzcOtwL9YBWbplWV3zrj1Vlzop05AI7Kh/T2cWXw
kLwDUcWBD2mmzsCkigjrYxatTiYJ6VvDVF8BIFwlxjRcvja7S2tX6ttjRNE0hcHZ
/hQMCIDmznGDi/o3AmofWn4x9T8awKdi3kYpOxTyAi243rd0Ojs0NCvHPQYUwida
tOx7RSjxnmiYrCt2bVl/4Le92Wgr1ccBMD0oS4oOJTqivGCvpNi0cIuAkmQEV7dk
vC7x7gv3iwqKboVz347Ju8MlNeqbl6Al416mM83bidy3io7bSVZ6BCUIkybxvQ7k
PcXP3m8gcwEdwaXlPmirOjqbzisFWTm1n0C80ljG1hytaaYfwqiOckIkMrxB2TYS
yO1IrIovHBxecTKUzK/KOhnsy39IqrYDdFxw8kEYbnHxZI4+pb8Lw1cRsOoX+BVh
pMKh5DwaSlBRKxhueuHOQt0LlnT62ngs2JNaT+zZBGZm9bv2sn4WPIJCKoZJ6Rrc
RHWf5zqYZ2uaOk8ui9OOJzafZgJbfORAF7qN27NsH9fTTk9FcsD111WSNTF5ANHQ
UBjPhhHTZhZib5e0Yd15dlZjITODN3fJzwVzKETmoJBONFIyYtl+BJYmjsFXgIlJ
zHKGIR3HVXLr/lbK04tVDcJHKAkOWzigmi7MEJZBd8/D1m3MvdGMoL6vcV6JVC/2
ssUK1lUya1xutDWglTyr2sOZ4oD2zOCBVM9YhPvN72fpM871ekYPMo3hKOVvtFYB
NCwkNj/QHSl37LprEjokSlIKZQ+bk+44Mt6xEKYVWDt8+ax6x7TZO0CLVE9WU2Nm
6c4WWt+kudv2KqDOZwoEUwzdkyEAQmzvpeHvtFfyXh8NZDq1lRkqi++0KASdSqwx
MrvCaBRupugUQut5gD53p+OChJkkqKuisgyB1Cm5zrTm2LmREszzCT0Pe5037Fcn
KnON53SOW02gBoe6nvWaPhm4T7Gov324+Iuv+JLkz7lxQvjsX6ZMyG8BQzpuu3ch
CLh//ei/Cb7f+//sUWT1oRsgUTdOUt9wYw9DW4ssyEjmc+D5RC79GwJFF07XB+jr
SYbKRag8CcVi8jU60D8gxNfODz+B8HRGAvnNL3xpQUJdc6QvPno2vTcltuuuQQW5
Nv7/9oIMqTL4gywOZXKSUPWoGSHZE13b2fg5ihS/Cl1WYBl0O+6QpLvGa6Z3jC8J
3QUUT+DWbX6tzx8Mv9Mcj9IOo4+dVfEckx2a/Inp/PBNi2oCasaUyBquBFdxN5g9
39UV86Y3PjwdIeFkD2IHnkvqXLDCv6zbNGNFihJHocQMv+fcW9qxdPDqroBDai16
ZLTlNjMAaFnxfkncHE3gmgTKzY6mU874X0Cn/4lQWW1myFQXhxx7P+FuNYQVPxPP
kwW6Y7X+5Y/dcYOBlAQBmWB5dD8oqXWHdUayL9/Sjuc/qCaa50XRSKgtRLG2l50o
zwK5j0L128LdMMXHmsiYfGAedY7AdCdSV/w3QjxsiDNkZ/V1ooDUEhCFtTfIjpcb
Xd0+UVH87pY6ERJOtAJYgiXdZsbuoJs+pwQajRlqcMkjeifOZDWihMB/Q9g2P/qi
jAix++II8uu+zw7U+1JI2YD41gqHbnfQd1PUHvvbi4xZusHuPgZBUUYj2k3jHBlg
L2vSOK9YhGfhIdvTujMmtOYpiAoHTcsAjYKJJcmmq6qLGKysCZhOE5HrUjv1H0pr
YyKbJzhaQrdLT03eEhUVdCzPlyBLvvwk6vs4b3eh4HgC1PvQBlwOAAcTOCwxYfTJ
5ml86PTEGIqwTsf8XL+1wzQpzIV7cebLrEpxF3KyoakOpVDSIhJcwAMuGLnioFDA
8eVVYlXlPBtywFQ1urnyv2TAkYWzkFHHpU09sNp0Qph1f9O/T+QNv4ThKu3Ns4+C
IB5Tm8DN0akj04zyEKG1RJhEgHaEsqPN9wK7Y+95rTdKjkaX1jOnZlB1C+Q6oEp4
l5w1cPJmkrN/IdR25CnEVzySNuHws4dzcX2mFyPg02wO2Top6gQUVpWcWNZohqx5
/ugEhoOZ0g0YcR7JxS4PUXRjsBI9S1O/t470jj1OfZE0nJJN25S8XYuhL7i7o7MH
wwhUMwqL9xLrvbHIq1GWzR9f0Q/M8KCZsMd0ZR8UfjbLUBYBn/+YB1t3xLz0YYtc
zweYSTGwX0L1hqij5Jcj5JCKXKKYXtZtGdZcDi2Pr6dFaUq3t0AmARtG77YAKC5n
vxa9J0W2xt29JlblTh95JnBVc3pQzhanMxCZKCJHKvhbZZgGmwwv0Yt3nKZnneQa
9YbwqCcIsDKD4b+RIsdwGR7nviGSwZgJx9QkiHxHTYq9L+lJKr0mMax9r6bJhAke
v1G+DOfK0UoR1FnisDNhxTeMdSRelQ4Q8gXFJO5UUpcE35sVtply9XYO8AagXHLR
mpJRWQTF65sey4WehMDtKAVlm49O2DbL21X4GvVtQ1wzAQVMdd71JjxxzMI7cQjf
mPDBZpGfvGnzof+8jCniKSaHc/6E+4ih6JDAG1lyvHhg7BbUgIpinKEwVHQ5p6Jx
g2HjHaFLhIGyD7YRkcCekHVWfy34yBx6SZVW78DS/qqeTASgNCHk8qYMNzRY4Isn
wIO2XQDOnmg+KCpGkVMRRvJaxikz8UCvwVyFHE/olaE0wpOZTfO67sUl3+ImoR26
S6m7FZ4jBnmS+OQ7qn+4EdXDPa2u4exLaeu/x/F+YCmV3s1aYNndovG2X7QyZSQP
sBPZhyqM2lpVulx8TTWzDtf9HVMRf2w3k0Q8+/hUsHPsgZkvWTPJUFaexDZrnxRF
LwIpFCq3Cdadf4wi+YOYonARdr22yGGCEkGxOvWUsZD0vVJNzb/t1rcMSKtyBgDL
/si8C7gew9PdChrarw8uVzkyITsUWIQqzUpZjSPWTHxhwl1CzlIhBHb6WJO5RjsH
rUkHLfLLK739XkS0D3sL+PtfsHgnkLw1vc3yIkaU+83Of7rYJqhjNwLKxs2hZ+Il
UVB6hgAWSDt7oYFU4JbhUGtekVKoanHhetSJvXqvYfL1440bpCMq2eH1GV3O5Ngk
3tCsA5/G8f87/jEk29FpAGqODxgkOVp6gB2cGvfICE8Dw3Ap7uV54Qtl2Y1tTKiY
9ISCsMtsO38C7ucuDwKsikTgoWV3PEKQzjMKbCBakDBYp+FFd41/IE8vEy6ulTiy
WFKQDEaop1uCXwZZoqGDQ4FxRavV3uL5JPaTI/zu8mNj2ih11SWOkQU7oox0X3te
UsUrz5gkYZA5bwQdLkWMRWaEdktJz7Chuud4nMoZhOBoS5wKOIn3R+Ew4iEO9vy0
9a+yixaTGOGhJPu6F4j95A8VMCcEydN9uEv9cnQ2/hc3/gH0iapOOz651uX2UM5+
ZGBW6SlHxuytzJeaOOJSV7T3q9wnS2AyhVxKED+qXaGdBZJdJhLJ/UxEQEc+d62U
3CizAdnx9cnb+41XVURQ8tVlKPRYz2kQ5Vkq3sa7Tyn0t2pzMu4EXIaIipobLFi7
Md5meyQrTsHS+mJyO6LNeqf7dFNyFa6qJATmRlIcSwW7Nl9A4KmKmWYnL+H1TZvG
gUdo26wEHLYFRFIVBzLL1fTtPCD+AqZeNVPkKKM+UXtl5Fdl/Q2MCthB1O6aZs/X
sNJIDIC9h/wwMwDk4M3xzvkC3bPabkmfuGijgJyeoxOUYvOhI+nkv1A++5GXVIwG
iRiPLVopZqUEeDAlNjKXO1qa4G/hK0Xij8RFEVpZ1ipmCKlb4luIOfoiSrEGBf32
65r7+W+/cgzbVURzsBqz/Fq4Vwq7aNYCr3UVUh3eV9QrvldI1kQzx72i8ju1k86q
xcVO8Ps9pAZeMhAphYxdC31JFhzgzcQjROeBsE50fOMpOKsGeW5UCxA3+Cm1O/zI
DQD0Axwhz2XrScT+pI69SpBdQXeBSNaBZKNBF7RtRb7mLcmX+0Kpt3x77jyw7DS9
V4lk0O0mI6MW76ljY3AhF4pFV7+gJePP20EMnLK+NxGmrjnswK6CGMBoLjCs6re3
DQ8EKHjCbCysdCJpxMehS7wepb4NmPk3LxAVlt7FQrVZ5eq2snqdkk4lc2LwgmSu
2PxT/IvneRj7JOjtsDQnsQRAvPk/3eKcGXr4ZT4bvXyANO98WFLkkv6f8xQp6ntH
RRIvooI5RTtxUm1isrDpMU8lmH6SNBWbFO1bCHFQZAoO09mQiLmFh/Obp5CGX+ce
WLHBaIUzuGxOot42JdzohmtiL7RQhl+NLDkIMnh8BVHoGk3saigAA+gldGxE0twG
3o7i4qKogL4SGejnsTZ9hFUjF8m25pu9KH6e2fWP6tO/RsxeD4311HpFfrHbCpko
Evr+sonXgb23nSPVqXi0BccKANWGc+P2u2u4Jr4b0R+RLk3WmYkscuo9iS1f1Bi8
GNraofw+wZdzslExtzLMJTKFQjgi+isvWojXuspdsfjGcwWWv/aWdYbafz5ZciIc
JHiB38i/DgEu0hiNzHpmbOz7wSLMb9akNknpe8211pJDYMpg4MHPnCyelvCoTFIj
LVBO5i/d2oAp1YXLUo9j5AG4TlhnOA1s/ypL9PGMGlcaRb/V3DRMTy3lZ8F6CyAh
5gDjX/hzSwPmXU/QLflxdq1cV5pa7MR6GZJqA84ntVNWmuJyjaIpVpawqQXV4U5G
/ENY9xgP2uVxUxfwwyD6IbqPc0/+7UaULw6cj3XZKfsDUlP3gd4JlSFlMuqv3VKY
dlZiS5MxvTtLpcYlen+Ab1GSl2TZ5asEPSg+n4z0K+RAjgYorcTAREqeZryXlTnK
AqySETrPc/rzHjVb+pPhGmf6xZKHUU7afDRVZEZz+u7lS6+fwPDWHZRYBEc1ppLc
LYXNpt0az7juxM3u9lWikb5WGVn9Umfb23LV71fqWlTjo+kf4v3CTWSSen+6pd2D
WvYWA5j6sc+L9zKzWuU3a6OZhS4wES6VW15YBkfSBZ635khUdjRzN16UUm/R6gNx
uwPJiH04tkmk0TevVbic0wxoMCK8/zj8uqDXFvynteiYZ9l6zo304nQudefiWjXt
UDhkz3rpc5RVFXBZPwhsQ1QKHxqsyjtSuebknyjpkgpnQxdxbYTOF0Fayo5J3K81
8TTb8M9MoX28jAkoeIn32So2opO8zkVF8lDkYTqzO/GfZHZXAYh4ONjsajK7Iq+7
w1E8btXcNXA4lXWREHlM+JoLncUpaRcLlmo/1S4eS8/t3cPc3HI/s1vvMwc4dEq5
SwnW3U9KV/qa5ulYUa/jZbj+rm4bymrWUspqqVolq5iu/yQ2PDB+F5rabdC5XS7y
6FgXyszWRYfXp07llByHlHJ78yxYbp7hxp3zYBdyW7u35lVtQiTKCrp4jveREHU+
5FLjeLG8AeNjrdNypAitjJAdBF3YxYz7RSRkmhkWsWqpKmUqlAOlkh/ZaUzpSkc2
Vhc+LwX4rZUDvOcmlSfFbUmMyg/Fw8YOad9YnuJOi/+4itj1IydRv3Njqd1F0eQV
oACy/YLUPUGboCBMbB4tYsRhDM87Rr3pBCpeHDUk90KEDAdwn7moG2tQq3AUdF0u
y2i2gwcfyR+HUdzqCyGyQ8j5cckViP0LNgFE0vRF05NyaOWdRbJVIpF7cpcei0v8
856AaGglphdVmtdtNVvtMCcBjjtq21Gr9I2UG2pyMDpuULTflqp9Dxr6WzBaFugh
Nm+iZ9EFgeFw8SW/qXvMdQKekVmXYmEZ+GbLDYYbWFyDtx0invtKl2p++xN5vSbg
zkbT6LXUJ9ig2Ms12UPL9UVoUsVXGflEMnhxvF75dqiE+KhR+n4ZTz6YyDO64f+/
8nH2/WKQR3vHlEh81Ox7/fVoRSebgfyac29oHMdjiYGeS6h3vxC9norURAXAqyo4
jKkI3BQq23VeG9I9i1sXWcoCNJahDCDsuzyELsuGCPKcHpr845ObPGhtdRhV5PM3
2V6LjCbMgvgmJYw4wSYPdWKtwZPDjGPq3p67T4f30xjOutaJ9yh4X0+MeGsoRiLN
Po/3WlODlAgwIjAQ3iBp/L7C6BwfuSoc9hP83W0dW0nvo0IZHuq3bRx4K/gxqOJY
xKvvPcxykuKr4tzMaQV7loS4BdSyk/dWQ62whUtWXfqG/rcEsxvoE2t+QFC287Pz
Q4I2m7VexOGyTttoEnf+ZTwZv7bc+9QO/I8Qj6Bh2Mp5QeJSA6MiCY/AXzsGCckf
vseXxjYY0GcpnqAPprkac9Pmexr5/MKY6BKN/HxA1gpItD5JEDTqBMFYGhlnvQMb
Z9yP9sMrslnXl4ucgTAw2MIVrMuKImBcpH+t9wKLkCB92xRziTo3BjO2G5f12yzc
GWUaRZG451dwLkqZl/48iJgI+tQzi7MsFNCU7+N9PXw+7N3O6JPpilKNgdnTlx/i
5+iMWB53sj7hqrQXlnVXQSXhoG04KDRP8kSZ0B1Jhqoak0BL+jpIuB/CkYQa3Kp1
e86lr32U9F/upCjko69+LINW5LcPT/YdcFQEAOe+8l9ybZFrPrmlPAt6+Anhzwo+
4jVG8lIKsSJcYsLNIP8HjZR5kiv/is/fjpUmOCVhOsg+VO67YUgxl9vN+7BvnxEr
S0GyVdhI+n/xTObNNhJ2TowbxZI5baiPXSzm6qRSUoHQh5MHtiWelpri1pkHtZQl
D+ElrEkvPyi0975zmd1hdhaAT5Pzu2cIfGGTuPFSMQIP4QAs1/JdFSYUAW1j+/ex
/ZEXggsqwOXJk3HVqoSyM5UehCRE0P9mMbEs6yEwuZooGe0XRSWLqIoyADSS2EDe
ppq3hSFqcoiPCCkRduRrMEHKC/x84SK7M4EHoQmW3eIZ+kYJKkQU3OLquiwDBvRI
5rKprKQCowVqPsfV3kJ7YZ17J88x9g6FSYMn0pMnChZaFrUe3KO06kzqx8TOPQP4
umP64MtevFkTgJ+dhn6ANBJo0kC+cQGQqZyyovjKh6c8Ax8nkGAmPHNtsr9k9iC8
Q0Fc+xENHiFcEE2X8v4G5ao74SDI6u8i+qQ7ak/Ey80bfCKTulL3OcaeZA2jgjEF
LMWQaKq3suyKbErydZ2wM7XORPHfFqNEEZY9Op1daiOciI/zxh5JkUZWpiWljRzE
NxZHj3nojJuun4NHqZ8BrVK6oH6wBUfyYJBbWnHuQh++00yHc0q7wQQbXMLYiwPj
B6+Rsn3NqJte6CeSG9/Mb/n8JaXPkbeXxhlXanz2vbNAnrs2VdNFMzse8FAsVWUd
Lm6XFlRkRsSJupnWwPBf3qer20qmrb6/sgr0Abtzyp0wdRkWhn9Bm8xrzEuXRYW5
ZGIWAY0wHNnX8uVIaahqECZxs7ILkX/hnpZ5eDLBGeIPOQa0IbtpzEXzrIFodx5Y
Iko3sYisOBnI3iHFIHbu/RA+n2tZwtyNUvYizN95tcW0uQyYRaUQCQtcesnFT4PZ
bi8O7RutxgLhf+gNeXfqvvAZjgu/Waun+4c+Osiss/AjoPM/QtAyTDDY+t73Fpuo
hNEfNnRh+HQoz39Q07e9+QGVWPKWPYXb5J1saCx6jk20HxkYpY0dLt1QAh/UsF45
H1EMwmMVBzBpjJxEflUlZ7hQpn86AojJ6Gv2JHK/HwurZVbauJ7WmreJDMZFkgmB
Dakj3cYN0TzOLCV60Hh5F6yxabWhyLKJrDmZ9LYwfQSyVlBbDKYtPElx7HRaalc7
XlKOTMAlIXs1wuGasAnVI1khaHWtuEqxiZgxXBXfuo8ZgiR9VWdQNHoijyIVSJwr
CkpF9ywkhm3KMgNd1PUyUAhxnVnT0A2liigvc0IihnCCgPNrlijEKic6YbI/x22N
cOjoaQ6yyrQ4G+el/NUxz9x9Nv1KRiUm7A8vA3iTNUGH07zOQAydNhk6Ys9wYNmW
zWd5Gu1+dM2Sq0SAFIyihAcyzePQMtwM4zcbMVuK6+m/xn+q2N7YwoK1IJrFFt/J
j/cPUzCiJEvG6zsGKgeRrqHGqTtW9q1rL6i8R0teKUaGZlwDtEfPPbLCpIkHZZMe
A5HSkDHAX3eyniR+ucKRZ/5KKm5yjMVxibSzsygli1oZS52fpP35Z9C2RITEfOQu
2AgdQBg/GbLtYoqAPgU6+MUDjO2LPgDomlaUZuH9Z+9EmT2Vrs0NKPwGnLXbbNkz
QDbcBS3ns7WuMmUGfRWTiLDeo5mTZxMVfLL1JgJObmXwNJ10zwfr96KHduJgqSaP
wxD9zTP3MVeF4ivIx2D7kUVX2toptPcxSQGE8pZSo1GZnYyehZkESIB1+s84cWbD
6Z/db9uDickJZAFpzVlXyeBz3AzATmVvkQWZAGR8KyRaHd2F071k5bHr6EmkRUVw
P79fPpBut5/Tv7p8xpjBTsYnxWUexbQOrZu2SqsBiuzyJxixM509xi/wK35upmB7
LINrf/7qNhvkYvX8SsqBOn/AZFpjbHC/pFt9aLhNULLUPQ6shgwAwcR5u/gDVGJh
AQaMDkVi2vxN/fFv+K3qZTOutiHGka+bYGsL4sNsizxQUpXm1EAj0IpQSNogi3wO
w6Zqq5gZsYx9g8RsPAgYwu8tB6lv3C4D3AnTMiq2XOvmqt9Hyw9iRngtQ/3IP5Ic
S6nPFwJCmAQpXEk50Qoy5yhuXxQpHijJxY0vEGS7eR7ziYHTNBKbRShOJLgjcQqg
+4Jun2vzpisvMoTnKLLDMOOGZ1COilLWFELj+8Yo6WfKEPCA0t5LTTgG4vbSD/Yb
vdrsSFcnDNYcr0vv/uLZRAC4nyRn2zNVVoj08fQml8TTl8G13VRIrl8Oa9zj/yx2
0BBaExqZOdHBh7v1L3YIrgKgmBsxY7p/Jdg77kXFTSm58VZXPaD5MMGdqDdC3oiH
t+HKg+nVOgYfEKA8eVbES82UhAGb6g3utLwuCwUeZROorUoQqtY+QcW+v8XhuGAN
T4+6TPVanq7ZmqeyGIeiHqPurilYxeW7PkM4OteHqRc6/H8xp64BDde2bNOcAw1u
PaiAJ7sXcm1Yiq91SjfbO95STavMtc7QrTyoB878YtFX8DdWPCn1jH7FF3ag3CrF
JRXUP6wrF9EKiE67wXdZE0Cd2RkAj6ExCyqLuzDo9tovHNQy/VA9mrcogNBO5/eb
qJ87Tli4rUSSKBouXleYA3731matobyFR3ABSq68/aEaAcMF0jUKiA8WXsJxzncN
l3/jSt87iyAg7NBVnIkYvRI3E0nQIQY0aQU2k6Nvq0YeAJqTBeDlSHMY/+tCjJbW
t7BrNb1gu/Mp2UiM5eE3t0bMjFaQE2bk5brtz5xbTmHNPGECQzuyAjXozy9MapbR
1x2taLJZKzCjVDUVaqjrEpB0MypIe1o0w8zmR51Uovw11Ns2OK0iJ6pqpbqQhTcR
eXyqPtviyc58e1HL9kZgxPe0syxGetzsx2qlo5uMtzA5um9ElSpS/O5EFVWgHHZa
XaPgbIgR5C3UL5M5ARUmrMQPEJOjgTxD6JdDMDrsFKfylvnQyIu+Cb+6kFupAdLJ
BmdZSOnq6fRxDCMjyGtNERqeLrJP7/TceD0imHaPOY8UO8KubV4/xXGef+V/1Hzq
jLYcTLheaX5LNDZIC5kJ3kXf5vM7RR/IS2OG7xodyA7q1psZlNQVtsCJi5dH0V0N
hb5P37EhmQO8hIXXMcbPxlO0R4mNpWWPeyO2H699E5IbSymPi+pDoVlUzSTnYUaZ
eNdsiP4rLhPbvEJ5OTXsUPMZBcoFgKeAV4ceTeya+U0ok/dcWANXVs2viQ2aCTvJ
oMTYmErBuL/mW8gSfc08+Kwu9KvB9YQaL8ulII1QfiVP65l7aEr9/dVFLWrQla9D
biMaWPFcirC/0zyfBsZdpi9yvgX40XY4tNq7NK7/YAYT/keIKAg0/9zaZ5Bf3lq5
4yvpq82CrIjh1KMmGgB9sMW+/EZ18FsKxypZRsiH5v+BDQ4XwRknorlD5ZNlZyW6
uDskUc7MMnuoYKG2H1JLzbMN4tVECdbNF/02Y1KRDpkGe9TVhmQSqc+9E12senfu
wrM95Ua4oaeF/ugUhYHGBHAqP9DXg+BArIkQwkVd7hmml+f1pX3iH/4huUNFzZSD
oXcE/Kkq0xjm1z28bTTHh26qKuyCsYdriKRXlutCVLJ4MNuu60l1S2QZyaXyJjoE
XuN3glGhpuOU7deWcivNVQkqLK/nX7nn0KiKESPwGQ7wFcgWHwG75xDSIal8Uqu+
HaCIqGepha7bh6hfDcqkQuEgHi5n1AjbHHUeL1HZASRwBsNFrBx74m22kacgNZ20
Rxeyf/RTKa+FQOBNNgfoN4InI9QB1Mp87Jdf4cCmaJeY3t1QYfT49eYzgD6RDpM+
7vL7kwallVICnROezzhNx/qIEpctC8Ua5SqTMoLchagUH8Ux7IiHL980WlM9y/u+
dw0vD/akDU4E7W7B1cTQATAbhZPmfqJ3kXwAAk8QvsMgosyjbdd3prNXo0rGji1V
bTpvK5kf33q41VwUL6fuPs5CiiIJfcghecvn0mC22YUxzOL2v9lF9/gMu7ttTJ4x
dXvpjpowCz+VTTOjLEP6Lm5PGDnDtcUmG5nub17lDzF3LTSv6lsz2HZavjILX9go
6VwfBPv4KMNL9otzLNsrRitnoqnFcQN+r/UsTg3ZcdIDRaqiP8Y/ETVFbnKQCV/R
+hgwfaELEOXJuwsmzMBgG54LICxm8NIdxLHLdRodZ3kjdgulSLkEWOkna7Kvc6vG
jqeIkcWRUEm++KcpIr5Vx0kI1G5xkbByjkedMsCygYf/KCLNOERSDMyTiPazfVTH
ZLiXo55pozjl9x6Cta4Rk8stsm314WSzPci+Dn7erTkaHDr0ywxAfTgqJmMkzeWa
egtVfhPQtVqIJQL8eiv+Y749IhjNa859+39JIDp83vDNCcd3spLdrFs2abUvYiDZ
wdfOshvWSxU6BN394QqeCZ2gt7+o/jCvLMjwhHCCR1l9nZoXYlS5CqCkV3/M1Bb5
rc17Pyx+mVBjsXyw48Z8J6DGzU23Olt65rA/7yhkj7NkrYuUR8d8dwjYZI7DM2Nm
XQKh8dBk6MiMljeqSeiohd4iHmldBhSEEDL79ozPjHpkKds9SAt/QCsJ8l5meU8b
Z5xoWDts0UjQMORrzD0sCCN0xQEh6d0Vvkqm9C14gJ8DSPUiAgrOf9XKOG6FslZU
uJh52QuaCVast2gfntcHsDagvFGTSMWmMo9Nip70fFvQv0z4bI4WSUG9kxOQfjT4
vaVzB7TYD6CyU0wQHm7X8d2bN2RCP/ylvyuZHaBxCtrhiDqEi/ljBPlgbZpUe3vv
Y8vTy/2p7M8IWx8CLAJz9aRz25/1B9FJrqs2CLhr1ql67uFmfys3pheZ3/6DDRxt
DB8C/yNZkf0ToG6yo6h2e+ULOjzCWy41FmEyeIZ9xsMz0jUZ/Db/opqXdn880hAQ
YKDsfYWK2YHPXCBGfhcE0XWs+Ted92bHYRUBx/jjPq5VLptXu0LbuQ4ctoMwleHo
AICvh4uVZnaNS6mErT9yH+YEFS6MnS4Tw5Pt0lZeBl68iT1e4L9MzuW7YZZDiSC2
zwyIAAiE8fy3vipbI1nnT3g1HUYyNOZaBeB58Cm3OxF81j7lrilbBCel5poq4oAg
7l+dQFh9+iAU4StT6ZaJ1CRKfvTAphtEMJmbtk7y7UMg6j7w8N1QbPOJlU/vyXFB
XNP2kGiF2DB9KqQahoBp/nDzs+QtOinvYLMkAR+B0dZ3E0n4PgZH5U3xiaTsPFBa
vCcsMQYlBdC3+x7dK5W/9nfRtBEaQXOInUEtDkJekxD4OhD6o1EZWhbieYAN6gH8
lFGsonYr/Etn5l++F675PNgsdtRzKui3xIKUL6CIC494LWtzK8zE06DUtUimIG1F
RGJgvPvvl8DzlZ2xMvLwa3y6Vs8G4otaHSavtnH69t8eZFFOk9cynsLfWZWyUOWj
hRpyCR94+JGftT5VyApUkAikjJ6PX4oYPJjz1IMUqaoODoe0GHQI/KzEtBCKsOBo
B/5SFO3plJRfMyR6pntjPoWMfracDvc3nToAYAqDXZyNoAO6gLLlucGd1amFB1GX
68cCPXpqPBHbFU4/I6JpJaH7s5m7p5hxNgcRM50UpxOFMKNEKTPPAJgAVSQ6QlQf
AECxlJ5VFq20drTEf7KXH+UAWtTq5M3cBAfUipNFj7jQquiKKQjLOmb8e7xOUN9P
euMWaRoR/EC7ojDDo6eNVk0g7ec6CWFg+3U77VKl+BlN+lPOR8+8k/JqfpNXQV83
5v4KGVioHJ68Uz8K/qf99N4CaXJz9a6qiStD2/vath8eao6wqZveTqY5f1j9QlYf
wj5HShTYrfx9aBbgotxQx11JXapUuCc/DU2lM9yNTobhi7oovXRGnAJ/wWeIIbVx
hNPyxWl29XZuiQlDLmMU5FcNfd0KKViEYV6Gc4KtF+4muQ+jGwNaCVv9wPAPFl/j
zTmOw2LYFYEgPkVJnLmhf6yBsdyjQK2C6jESmMonEysBylNrPygCnI8mPr/AeJMI
futt1GNhyggCnbxZObMtovJKwsbQegsJRWWDMNr9KWMD5iXUoFyW80B9rTTu04ko
A1/QV2qfC96zT279WJVp4lNt/l2VYlMj+IsnjxZpRFelpzcFk7X5K2WEnLuuQoAe
J1PuIuDEPY30e3LL994Spp9Gg3Q6n6TXFeIjy50ieUJLyrX/qjK2KlpZk0Fn4MSf
5hkhKIHhMyByjGKIe2MWg9IFbL4apCTvfByhIK/qetU2Bl3R3c899b8j7/7k3q8b
+iTmUrX5qaHh3p2ndVgsyLR23YEEXfwTKeE1gAdBK/YgRqoJbOzYh88ni5KWqwWJ
oztbX0WsTPDynIE7UP7cG3pB34iPrUzTgIZJU93PqbAbmq7ZnJFV7jgVh5qVxYN1
7Dz3E1X0gcE1RHlfqza+iUKSAjL1lzCkbwmhkKEkccePFldvuCwtXg+85lJLSqHl
epr+a23VWB2iEAf+IJe3aF99jcRw84dpB9HEcb6MOphLqRBihjAgdz6hdju9TvKn
HE1nb2OwlQM9P9PmHAFz6R3j/OJUXESPdrzhI7sRQ8QymeD3QbckU6HUIOzv72gw
q4Scbg7MEstCkXH4kiMz/5nCNHEstVxGkEXcvvtIDAOOlr7CsQCdQuhLoWYPR7Ue
x34rjv8IlPz0iqicG1qjkvfsF/QPPuF2dT3genJtdj54941KQ3ZY8qHczgc0Uarb
y0+B4b45jwA6+epUXyPL6XihxG2DDKuvR51vKVRMdEalXfRp0xtePDDewKcknxf5
G2J1ZGPjscSj+ISzVQ4dJRcBcfo1cLTJ7duMKACnVK8oyx3VitwEv5tW/gifiQJ2
vbymo3WZtxu+EWgFBP3cbCTBr6eFnRowdtBPO61lrqPZ2OMVL0h2NRc77D1yctYf
Xbo9Z/vnW/8EZ2356KwoxJEPNX32UCBrVS/3vLVT8DVX2nNLzzy7oohJuBIFkSNS
DfyoYN1nH+dV/pH0Jg2nryDECPRHwqB026oTkk5BMiU0lt5OYUHCfy931JOyd7Md
WaQGz0mq0032Ylo9wA3V2pcnDlXTzMyQjwnh1qDKfKSamlBCPDWJ9xLUqyPGZPur
kKdkQewslkZ1TyVi98TThJtCND5PAvtVe18fUBzPGTA7j+Nt7Fy2rLa1z8cxsp37
T5jlVzptPVgh3zEq26UXFiN2XA77JWK5fS4/BGLJSBM5u2Q07hS2Yxdx+vQ4ZZtc
sJc93RR4BCora/UvF2QYmbUjNnE7j8uJF8jL3niClEb3YMdA48Obwx4trISpS5w1
7KaxQTj0rwyhHX0r+027AZrVcaJY0QMmyi9R9+l+olLJJ7CopH/wSRyKFhnGeI2S
V5DH0q/J3oz1SZ4kwu82mTxOFfN9Ich6Rpc4XzYkAsaJmR9i3VnMy3gX9KurEJxw
fGcLeQxJC/Pv7pU5xyjZsVY9kMLskumEin6Y1OCr5CuPNHStjJJyobz+ER0SRT99
qaSaT7cB3Z0dUNPPe3XT1uj3hvYgk5E9nEwVg8cbmBAt+c3Y9VvqytLAQ3Y1iZ4C
VfOTl7sBYtRIZ6rhWE1Z+sA2zTXL3oE9GtXwzaPDZ936xec963dBbiALSL0HQppR
y4DKjHuqd6HDNKxJBXsyxLXVeFfHH3zE65JqIeYnM7zZrav70+sfXkyGvYHWTYh+
bqv8ynbZShrseQzMlB8wC/JI5smzxHZb0bAiRS2G0yB+B7cvDRcjgO4AXNuNbzlj
X8a4OQXX6DfTsmzmwI/vXsA+kM+Wy4KlGo7zwsQ50T61H5O/vls99boJrb+7NWBr
LmTIZ+KOknmCu0WppZU9h0XtW8vQ9c8ai11YkJ26yKmbIA3MP5Ah9d0s1YezrSeT
/7Bp+Ba9K/s3xUGim2LoFjcUW+ygbWwISwfa0OD48KHXTrCpD6971N0ikq0tuaDf
WkJpZaZP3RaTrAKWRYWmHgB7+cXmCA92vSbH0c7Y7f+iDVESTHecg8CdIuVQwBvN
dtO39J7AHJezKBsq0YMjIRnmMBqG8AgUwERqtyjoGZ7B3rRwcnKFOnou813w3jz3
BazLuT3WXvu7RRaul3JT9r5l9wEahFw703EcQAyEs6ytGnJh4x+pquQ8/f/DgScU
zZq+5RJmKAew390CFjfara18d8ZnvPykR+b+CS1DjQGgAnyA/uAg4h7GghR4AhWJ
bpMk+ddfZBfnXhcQl0NCpc5V6gJPJZWJXKbGFyJp4uw7IbJfGW8wQG2JiGUraJBB
/hflCbYKSbH/MpV9qy6vKFzNWoA1YsBqHFrO2Gcs3Win/wukntSxqDvWJNf94fSC
ESUJ4wUqt55hMbSCnMCAEPYHUwsJ7Afh2mf/5hZ9hIJlv6BY7SxD3GYqTrYugVgx
mkvYwm/V0zaMxXWExJWqikWZ557kSYMVBQ4Bn0+jtvRv6BcKSae578D+cn5/NhDx
k3SmY86pTY46m6nVzVU36l5eh6QQ3NYtUcpr+oNFAQ1Pje6PfW26jfF/vgNzF0Sk
sDS8Ro5jtEFsQAeIa22g+EKpB6iUEB/qfdvk7LRUszJRFmo4FuBjAY9jE67Q2/57
9opzAOgWfu5b0OxKLLez32S4E+JxZk6EYZzVvY7sFpkohiYzviO5AAFh/z0hwdK7
zjk++8G9UYmqlTbDPAqVu+YNeRyNpDuBRRWtFi4FnuokGPuV64cf0UJQxfgq/N4F
HGv+Ppv6fmhN9g91IOUfmdIavBDowtNycY3X9DJxiLs0MKJcRAOozEG8QJrY2A5G
+v3XN7a49/9dXDRTU2Fb25MLwoRLKyot3c/sxh0rbguu39LVUeQQn13eFVjL/nXk
NyggD2eHHCMUTnPP8xGf8OngkzygE+l+vaRqo/Nd33ufpi6hg9rCd7uGqu6GfULU
E2ODpObTU7JFJBmsAIW9cWtGv/SnmVDTRPaZWFZceemN4WmlNGS/ZWS2Aa9BtuU0
xn+v21TEZxx6DG/Z2Ji2dxyJafqOnyVTcUGj1YG0ThVIBs1pwOLlpoAaFaocgFuA
mlsxV158bozO/PUIuc6iJyigZBu/BBHcXaEVk/bGwSV1Cyik2118einKEUnCI+8v
57W1laCoCry1CUj46tPhFCiNnj521B0/d6UCYR3JIqeE50dWSp30pqql08xX64hY
WOZcmS4k4CMUSMBHQeZc/THrO1qUolsdUlOqeV8V6dmhJJwlcAl7kP65oWypfzsQ
iYZQdoKXZ9p5cC45cf29RlBKGEOhkGYbeEp8cSgPK91wMdp4oMs19S1inVc2KW8j
1ssQZGQch8cc5ZleokHlCG6QCebgxmuj+OpCiVQghZdSrQxTxi1IiAryEKrH3jwf
IdF1I2ddhgK0BWMWIEkm189OuLumj9hW4wq0lA1erqycP6YykSNJcTPzGshv+01g
vOfMylDD3WIk8H0zTGrLGPdi5M0xrgX4+JaDmGcH4cOrQlpCQR7XLhiNxJ3pwgyB
hnjn9nrq7YUE8SBhW6oxf42tZBrSVIvvRWrC0JUQ7GXO3pUWagKh+2d42odNf9Js
qEMDwu6zr5SUZ//JzfETRU8FKLq6xb0rHC0awuYW9aTs+/tyW387XpYRtm9YOF9X
Ey4R0+cb2AOcP6ljO0lmRpbTRpfUtcnTv+CPrp+2ich6h/ni65nMCdm/VY5KK7XS
F46EbMEAPvvGvOKCJIeALIcUAX1615K3vm0QcGXYVcU6f6m4EVxl2O4X6HnCIJ4/
TlGsBCbED4IA5NnUwNepj6cZcYLsmpSaTKJrnWNafTn89B09O/UTLlR5pDTQvYqB
WjjyzdRAyNQZntVbimRs1CAoLIkrv7MVMMwMol7EtWRzHcJC4Nk4D4JRNiN6QM3C
tQpmJNjTKovNspmRnEpUsFVFx2xMU+LIBokedGrYdRzoott3tBhT43prFgQncohh
u3vS9EGvRhrGWzM4BvEbd2w1hDp8tSIDHnJItZzPp+UrfjY8ZVfRKxa6WtrIj/O3
NVWp5p/J/8Z2J6rtKOP/hH75JjngdL2MQauvbUzNq/e3J64kqOPjVVuXh1B7EI0K
6zUkVCja8RPy62uhMDeXl+Iq4b4p3iFLC9Ob8Ur/XUi3wnenJ8tD0tRN5EbVIixQ
8LoqT3eKNo6jvUEhjWc/tLAtQyz7ARnmqxngC5Rb0hg2v/SCWqSNpKtu5IXQhBI8
uEELA8OTvrkqPc3By0OrKpAiQR/4sIQWpke2uOWptbXmd7mz/d3U00Tz3NY6LjeR
/vufq/leq3ZFmwdl69EU80ylO2aHp2TIOcUhvva6TBXRVhO+L7OE9SUarlXMJs37
vU9zZNlIkn33w5whZlMXuCxRSfbl9iGhr05sQv+MZewiszTzdxU1pM45uAeXILQM
El8dW3UDv3k0/1lsjY5VxGZg2hAE9pBBkG/K0H1JAl0XsqA25PV4CPL5fWfGOzwK
76ZjNMJ5EzdqS5KtiOW4GGeg4Vf1vL0FpfO6fNEmJvzs90BC7GnfgOEN9BOMtKHx
PcTkCVpFoqU4rpOZyOcAqQwD6AJTGfHzMh3RcIEQsAVT9vpA5FxxDEcFpbZ5hgRW
9M2iNisDvVc2O46vDIIK0LtskYBM0mdZW3jvu0m1W5AE1slWXQg8liSn9DRKnWlO
gLBHMh9GqhiJ6Y6bl4hKDiI1XGdYFjoEYXiVrc4XHc9Ny6cAxv7B6rxb7ez4oW32
NDOHu77R2XtGh3z2hBYTijtpUlQ2/T4B5x0Agpn6xuUOMHPKDai5C6SlnYA1NY3j
9YjoGmUI1kMVRn9Viofc7Ee8gzDBzfx17hsDJ7RvcEs/P79k70GEMuHhuMoz2Qqa
HgEzhckyHslnpeXAE/UkQ/oRC5wyDYmtOA2wQk2WjWeM8YCvwk0omyub5Hcc7toY
pr+hSU6mHoLa2n2DpMowKZyfYRtBlQlD5DhcHZYJnkvHw+3pPcenboXA9ZCi6uI9
uFUmKNBSFtBGEh4+wHm9So8UT0BiXTIMSDV7hft3hK5HQOOBCAoaw6U5QWh4CUh1
bG//VgByGAapE/FGeeDPm1yDWDzS9oQxDwOqdXnLJCsPpycyvDFGR03CRIQD+ONK
0RMAfNc1X9d/qzJ8iGDdK3urA0QfBg/kYQMHaau1zuiLUsc25RHa4MxwSqoQqKK3
igHBSSM5lIqN1evgeonM6oCJrl2p0uUgTp5Itvfl3oC+NS2EqjseOW+eoIHUnLxv
jyBPtKcy4KhtPgGkM6Gd3FE+3WDCL7S5czhIgyjNzEfA+KYGe1zp3R0JWJ+hOUWT
W0iLg77jZpb2WLkqHHEEFzTZOecYp4UNmiAxlK1O4ca2plG703R4ZMsyuWvGQjkk
QXl/Fkqfj/a94+WmWLLuZnQPFfyTJXqyebbcp/W5ca+n9mXEpOib13iR+XVHwYG/
Pq3TBVZuFRXvvyPmnwxc/iWFxpjiodSiL+uvYBFtOJU8fg4sSdBm0OeFisscqI35
EICbZ3PB2+hzMa5z91qVlUONjsMAdy7ad08LDoP4JZG7+gx+5yOSGov2UCz5i0OM
Ub9ik0bSaC3ZyFokOE1wiqD17GF0nkHtstL7jDcnle5iiC0wuhWOq+QOJdqJ7sIQ
9BgCvUtxMZ6kqJISAYdpN0AmyO9bcjyvc8qjrqWcqOhj1xUFHAHkiKasRzkHSyez
DFy9787WiiPHuF3DOCASkXblJImd5H2TyEIWecVKVU/v8A45rfzR8HRYBIE/YUx+
NaiBhK2SzOtOf7j+QbHXyaMB/VFWZkRozjZ0zgZ7oA5e6jhSo/hI+g0mvnK+xCAY
e/G72lG1VYmUyLdOGItYFAcOFcetE2ztF4ftORI5qIOaigFQt0d3fC88n1NrUzfm
TqWVeujoKOBBUIYt6zHyYStAR7PP9czrPAfO6Ux+5SaL4ppMLANH0QxotngtHGXd
UUTL44LwE1jdBtvtDQrvvFhGLDGreXAytzwwa1qUYy4jImIAsZvZTPw8Bp009upy
E5RW4Oh8VicqP0ybbn0bkd2J6qXgn2gHibU3JcWpyR3JoYPwrReA8GES0p+7U6VP
4qu0kGlWq9qJV2qXWZbUSf+Swvneat1e5FDoXqeCXkBCIGYODo3D3WMy9ZzFiwws
94/qqFn2bRUFsEB9lr5aGVoZs0PbUJ76tmSY3nnl5VeYMBBIFYUIs/IldHug8gp9
c+B5+D2T0Gz7CjJjny1zqe9TcNii0pDVAe8G3krmDrk/K3Y6snm97f8KqTH3bExy
9V/VbpPwUbDg4pbJ3Ba9dp/1SGWY4VBGXHGXWnIgljEycnNKnxR6rndpM5VgpEI8
+33iODW/6hqtt4rr7ERNOr8VXTpbXf7rKbjbSszjZtsSWnYbDTxyydylBkUMlqdM
YifQKm/cJ8EqZNhyNNLpGGQVFTPZBQ5Q3Qp7Vb5dil53ijJAJsTPVBu/1Kn2x15W
kko0OaXPIa5uk+QzLppoy64AvN33rcJ0cIzSUUWuem8gFXQ3B2r9ATToB/q+oEkv
EsMug9C443s4mkIW5blTXEJeyzx9/tdeFmw+PeGi0xQw9Rr7aybxHERenpsAnv9n
+F3jiphF/s7g8Y9p8BSWUkPPW7vYxCIcDEFKev17N0rSo/s3If3v9lWNgq+Y3qSz
n5qlYS64HqhLvpz4xAfe9kUN67u+7LnY95U7w2Q/KOSNFLmCgmIEBUxrp9GbmhqF
+t5+GMir5KN5zWxqGBPbtAXrSElqejzCnLOBl7lRayOYzLCUMvMHMfEqa64KndxD
B1OPwBfa5H9APXywbs7AMhmrIgKQBWIxFJQ6eVzXOpmszrmMdj3/ghOkqTEroYVo
4iKhUuTFfX2DnoyxYRRD0ptTWGLrnpmJDlswBc7u2pTB0orokY3JCLysJ+bj6i8i
CXce2Vzce6YJAz4DjLezZcs2U60yPcAhLT5VyDRk2KwQ7hC06366IFCE1/Dbo6NC
+D4ujUW3CSm0sKfJpqf1qtW5PGr1uqgawlZczR+IM+w7C7NboowVYiDPHOw6W/J9
YovRw2eYGBYMErKSIMoCophJlEVD2RpwGQivQIlDA/EvRX++omzQtAawCsW4Zz78
EMrHlIrHPcoNdDli4tQUBNnCKqA6/U2zO22GhEdcQQRW3DfXY9xhDpzMm5lo7TE9
cAY0rpKnUDKntHeisSZwFJ9xvMTscA5Me2jLGfW+vx2fzbFbidCD7iorir6xuMeU
uZxCO4ZPlo5DpoRZS6Welfo95AAsr3io0nobzGAUSP418Z/0GWFrWHG46R0gk9so
9CmhG84qnO/cvlhXYvL8s0IXZvW/gYAqsYOVWwmeKyG1FBLTu+QhSEilJunrY5Er
nLJ4CVN9bxnZ8mo5YYuLZKoZlF6wKZmyxwnpd/Qnfnpq4UImb0F7G814ItgrNafD
rsWrDn/KnSGqff0LXpOVbEyxRKaU5LJhXJa4YCQOZMc7yj+h5s47cCnWyu7I/NJu
U6hKJmMle/Inc8Vfn6uIheBF+e4oeEw6j8nScNZ5bVpUGkhkeO5KHe8TA+0aHKf1
dMO5XVCgTvdNHLY8asL4zVbc1yfMIc/YLCWzuUr4uBTMbY1zu94DIjXH96f/6Y4z
k/aKHB900Rate++RQatgEKc3ivrJu6l3CHl8mn568WV8Zd2yOCMdbvgspY+43TR7
+EBAnNqp4Z7TO33qjQTaz/kSHSH2oaVVyVyLby4aK/VtXfiJUrKMajdIVRXRGB5o
fjzanVPJMa8eOvG0Yt8CgyZUzTJzFd7IE9IWx1/lGE+daa26a5bvKB4EA4gkR2+U
kTysfyXeItG2CNnfXkMTslltqSCCVxPJ0dPFeDfgqm53VAIRe3SRJZ+MhDKx3XZ7
A7tez4eo7XwwQMImhFlaqaHhAvS4It2WJJExdBfwVbxeDhxBiIMLOKToCE2LECJP
po9L+cledRxi86KRmj5K+RlpNpmoINMhV/8vw3B+c5j6iiRO55SMRaePADbZll9Q
rn6Qw+v4SVYAOCCLZfWQTNFnPLoXd4XzurDaaiMK6NVssdIJYNfEcy0qavdHXWDa
ewlXg8dnKzdVrAQrS+zub5PEvhaJIwkuvVQeY+uStg85ZMF/dhUq0eBfY8f/WkkZ
XU3aytfrxXSEkp+zT8e/tjFEaldIvpW2eXVS5y+bdLq8K4HaM3iaYlP3xLybF5Dg
pYGKy4YqrJACmV4aHw5Dgr4ZiCPqr3xlzRe/WBUeQWfASAv00PiTCLVuo0pnl6hi
fnSJdTaGWAOhIIId5VOySnjjm+qvMlMsC0RgavofXEfHu5DrLi2BJEcKZWgqmIzD
A7Vps5z2kqZtMyMascZ0NVcTKdMWGlEt1Sx3eQGRklaYgVp1/Ukdta3nPedFyRXc
0sFZmAUGCrGOwYnsKat41YUXjF5Cy7Vy0KcVYnSAr3IFelb2fGOBav98ropbt8nr
wrkx1eoe1B1HXBBDeKdqUoQ8rQFyOve6PA5duc3EPCppG3WuAkmEPQU2QyG5ApUr
M+SeTYTxNAHefcU33a1nKpRSxonNBCDGJ/hSV7NdGP2di7eHz4gNr51BJX+8lYty
+wyZl3wVMA2hCtAeYeWYlVuw0hV1Pj9aMInde6U7GiAr6r/RILMMJbfAjL8XodZ9
cHholw5yUn+QGrXLuMEG22y8wSM+XN2OtQ5zMAIjuTpbUGv9Jgey+3elYdcUUgZu
b2OKZ6b6WiHYXjonL175btEjTDURE1CvcAfOwv3FekKrRlWcmaObxHkiMLzkGnG/
YyJlbfi70Wcpa8h8ogCe6PfWR7MGUAeZBWG55YSQXVnpNRPl4JGAv8Fn5590dVbj
JAKXk8EH3aQa2agZZyy+jIYqYRTy7s7subUnkYrzD0Fr2i1/sL2AgtFKWv4qRfIQ
OCH8B9QQczGvEY48XtaLFTxb3VRe0bjc4tmc0ou8dpXLeqW3qm/eG6Yhuij0evRU
w9tPzpcdE0wk+PkGrIfwPqvxHtj+rzGs7QgGKZfpPMf/jMZXaWwFhIeKvy7QgabM
S2Sr0lfoQx4aadVsPgeVlMf7x4YmhPhH7L30IpjqKdLgU41YQJk+LHrJYWYrDvZn
D2/CSGaF5316YV5Qq3aBdaTKgElTOx/yiSRhqyHebYBV8DEbiZqYBtOWSk0ADO6j
oNRVfKdRb4bcJXwdRJbdneLzjmXR5K6Aym71LxWgtcEu3gSgvM0nWMpuMSSeAx9/
l8RMUfOlUDHeClAM70qgrop9qng+ZbD6ACpIe12izHOMEDLmQzW+aijE1gDcCfmA
vA27/kxwhsKohjJ1JcoDmiJkICMU5w0poBx8z8athGpIresl6BwbAf4ogmBXBxpO
e7aaTqP1lBeDn1rwxozmqKSQEuFfGDexfy+KFNrCjd+lMFpwFygX2cgn2ZM6WSmm
UUIv3JKFQsROUT4aAi03phWUMORJhWIIgwWwDvkbRaOEhxqdTyQstJ6Yl1IemP9k
kgj3ZqJ4RaVjBwcndy1uL2Dbcz9cIAcdVSEcIhd5YZWopOstxnBGeyBnxtA5E/Dp
NUouka1VYLoyhF4LsxOfoFrW0uESo4G8NbA3zz7+w3Q9hMaikIOCgqj5OHyRZ4+W
ccOO8RYbECiPYchBHuFnDWUXc6qwLmHuDn01bGsMlERueSSxZuljbTLBGKCprQ85
F1cK2RS5kS3RaYKh971kK7VqAdagmMUQKl6sfIYJN4pQfc2HX83620B8x+jF1M1v
r9+xjCrx/RL631tBa31By3DnHStC13X6BVh+mgMakeTMnZamkubuKNXg1aE61K35
EQZsFqimQnAgsOEvMiRUSenGPxdcKVNfw5Sm1X1fUJ2FSryhj+XVq76ZY/YK/7Fu
raj847HxRrXb+WZeZ7Qx3QaOhSME8nDGevijFBRqqVCn0xX17yyDkSjxqNuP26dW
xX9v/CQ56xD3R1W5i7yjvRF1P15lm2iXV6rzKq8gjHiadtSON/1qPm+kV7QpD0XD
lNDTvLrN87Yc9YIEAW5LBnRzNGafIC+DJGnONQNUGFf/VN5g2hTN47Gy3YgTtE5X
8qfppGseqRK5nW1bfqiegu2pt/0ZYqxxtoHr6Zz/4xSFNkOAAi+Is05WVQxmbZCk
LY5BIWdSUL7/yjR8ebXKK0OMvFmPlsk+hFeHZ/zuGapnpbYz2GqwZ4qwuUVSpWMn
lfFBeQNoQz6psFUY/hihNwXpTiPwG/d0ByAF/yyqmsF0/y/tN1oM+8136UaMFDWh
C/qEPTMlfPEYTI5dOZkeJIEg4rYPROlGcbxLjd+9tjORKABTqDbLPOu1ZhK7aFKl
xvCfYJWexnzy5C/RMxJut+9v21A3iNckfTr0Ql9+bh09M2hj2jNP+0HA/jBiGVjy
3EPNjneRdL65sDgp3+EZ4UrvwQnLrZYIl7dNPoIEVSHS+NwA0771kmKBGAs3acT5
nzIjqqgV02L7u/V5xcgoRjF2XeVHHBu6IFLOFBmWYoFhHI15H8vvPavWK5GEV3f3
K06JRZxZb1FU5eu+FoGXTegpJrZOW5ymjNXloGOWXu/OJOwM+GtgD62f/h4hrtdS
330i8tYY+ar2tvW5u7vKNH/Yc2Oa4Mhz/LLuo36jpzGZR1q3RgXN02L90hBC+9LF
vJWefPUPC8/dKVZy5383e+KisgpJFcotfGs1WDHFCgUJeWeSUj5RpLzCpRfvjKje
zM3mrMWnOi+008tX3MS8xOQf7cxvLMabvzBYiHgLNxI9jE3WtIK36v3FvsSwp8Tk
Z9KS1aOaes8jSqPtwWrzqnYX6GgsskhU4Yxni0YNczqv1Ivl6AYrlIH1qH58226W
YjdNx+qHj436wR+WAK6v5kcRf5BPDJqI8vGyo8xhDGAiOhXTWZwNGGxEqDUuxoho
zIMD1XtgsCKlHrD0Bl3D2M2AT+ThGygYjiWS3RZCyPAZOpqTyRlSUZ11koVIvmn6
EBYMR3vcuXPHHaA0ySNXLO6uMXf7S4BF/qDgofEmDJT3f4/nQAd7hwek7bct+0Wn
w0ACKf3gNWeaZFEGzOLMLzUNH/V0tXdK1IAltvbU9KJDTFlD2R2nOkexrlpi4FfJ
kyPI6zSfQzYf3/u2DcEzYPtxSwNV4KRqNiEnXY36S6md7S64u9N+EqhjdMC4Hmmp
XR8JW/vD6bleH6cfpmOAfiiauaCmuaUtBqU2yX2ety1NeAqu07FttM79GQhv31pr
QnlG3avCdJTn1D64DX1NgQZOZxIIr4dUcFYKOfPt4P64vFrA+pBrljxGBCLM+6RN
KA6W1HBH9Kn4SXRhBX9wy0db/6lahYeVQiIysdjtue+Kulhtb+przffYEYWj9rIA
F0ayr2oJETenG7kc5j8ohJofGSE4ncOVkVi3jEHHP6oz7WUPVMVn4nptR/Zggz+y
z4h4GYF6AwEOAWidrN0hrO8nY0mZctLXo34ABgpgH5ZjSER9MLgwDXO6dWcoWQTh
5K9RBTHb1MR9LfKkfFP0apjgCGAM8DLCJP7/W4ZuKUDgLRmNeG/oiD/7VN7d+Y93
BS+nCVv2ClWh5rGmdO6hd19LiB3Ku3dIFhYKBxTc5gwimGCljrpBgLu5WH3H/GD3
YTB02Bq7qAc3PDVlm7A+ZQW2au5nT1Tn56XdAmUuD1zsU9C3AhSDsCTf8/18qzAk
SAO5DIsFEnEfgCuyshNP3k0dwfGA98cXdIybdAm7AzrQh7LLzVLLsU/6PiE57RGE
RfODfNZ/AJ0bYzsiX2VBMgzpLx+4hrnCBX/A4gMWxtRt0FKLExyWd6mY7E+IuoxG
0YeYzrzQ3wCeA5ySeSxX8b9Zb3MwIkZMg2hRz6Vuy1GWMwclFA/T3//3wbGGmyBU
YAeWO3EJqWTcEcOiWC75g2OzxS4i92/XBZugP46CeyyEXYs+cShl/yj1geqRJE3y
eoEMVklZwQ4foZsbyf0gw/YvusKBkacf8q68te1LvW9HSZcqVHxpJi8kBmX8WKyX
XAEhyOl9e7adrFprasoFyU2GjcO22Dk63T07RAse2Xz2lFMBboj5B9UewsoYujnj
UbFL3Yj1fW1xxpU7RQ9jLfHdCMfKW4gIdW3RLcTPBgg2pawTK09hIzniUMOcJjVb
JRqyF85zgGeh3PlA/zKvntQrIYQIQ3CDRLb8e36Nc9EbV5PFwrg2YmOoeTbLo18B
p4E0rQSXUVCY2Oc4pL56L0cA7LpjRqmoCz4zccoDFU3mMz0UJKBRylaYXkpuehuX
oQAgNQIupvLFfTopXy87GNMjM1U82+2Bt1cO3eC7Srkltn3sdESgl5o25C2Z0ZM4
KwmmFjWH2v7FLxqImIj1gUuwoYvLi6TzyMdvOiuUaUCXCuALHpovNIgzPLXqBmA9
nwYOsbnDoJMfbHraOZAPbicdJQrZ2uup/IeqX4X5P7YuOKG3/04HHzL2Iabmi7H0
eyQtrSqeR1txkBB4OpZPDZITCQA3Hv53YhN3cMUtXFrGGeXvLsLyUduO5nKpGmPH
Kaz+KKEukv93S6GhFp+tBVqQkQPvt2oDBpc1QdbxxPeD3DQbD6b6wFFyuRzkB2Ah
gcqty2fPfnZYxZ6nqCFx37jFgHHzhADUPpgKMc/oLx1vHAkRoNDOV2T1Cy+xF4KW
8kvTk8R29QwSZaqlWrGFO8yf3gQl0v1vh8owXmRk2qFAvxZwj4TcSZ27r+gNoyBq
5qP4STLxCyXG4XNZPUXKDIpPLKyMoeO/Xp+VPL4MHetGdlHD+Pza1o1CcNgg4D/t
mOdB3H53B1R36OVQKS+y6HeaYooDtcXGogNjHCzUg5AFYJAXEAXofbtmguUke8Nd
6KAtYqx87vjrvw/x6S71ICLBsJ6Ua+TLSDLYx7nqVLYmu0a7HYZrCwTeVwcvtTQU
fJLrX54QUaGgEa4l29GSZGjuUldf4nlLbAfkZrcqv6Ab5s5qu/VF8oKn+M/Eqz+U
rhh2EdKwuI6HzvoSQKHXUkxx7U1bNhkJWP/Oi/gM6vOyPSCJ1+EPJSvgvdZ7vlYs
MQioBYUW6GlvflvaSJPpVt3TKwsuOmvSf8SIMAY1SyF7/Dadyd9HV3RyHnsrs17x
taANO7YsxrmPEJ43fZzgPIKBgFjRtLaZCKQzKPzqU6QyRDSLvLKz/P7kL0HSrBN+
9FYgXMOAIigKG1IZbiaUfW3I3lvKOJYIc6oBX5Vr2g4/9au78CeyfsK45vDx3KPw
2phRSFHjDqQcmeoWRQMDMt7pd8G/Kp3n9c3AcLZeKDfMldjSDYe0+SzR0TE6JSnL
3Ta23qZ3DAziQJIiTvDRRaea9eyOc9Gq50ewHzZ1HH4OmeAh/DaQfLh0dAsbQEwb
mS2SppJL+6ECjNvWyUf31IkGJ7UTN5U5m5dGrp9sbhzY48yOlJT/JzJM0Lli9RaL
QFZNIjkRvUzCX0hzEwW91N0jW5MZoWQURUt5+o/rdeihAvtqSWv3NyvPSN+ztzhq
uNKHziIBxHlRuxzhT7L67EEjPuQrQ6uBklP7mFMdbj8Ntfi0Gmj3W5Z8EoY0dCzJ
4q9qakty60qns2DB1RAmBeDzwo28FFQ33QVbNkJVaB4EdEDScpdtbO/CpUWEifUx
2Ia4HQc8wvnt6VLARWJmku6fTP+lJ0om3B5aNZuEZ5tZ0St/XK14/WZ1T8JvvG4P
1giQ6Aoh4ZYk9vO2e7ed8sNHcM/30RAgnTypirbcZYtetwVHLQ/metd495XC7ccv
48LT3zFHVESH4Ih7BkK6RtG/TEYmtHT5lfrIKl9DDqSBqWjzzW0/njMPLoqNnNxa
tvkaxDie81W2dNwS21Gi9KUiFjslzYfZXcOchqjPB0d9ppnixfTQCd6lGFSWnJ89
dRKXyv1F1t+x7+D5E5d9CyZ5qxhoITxKgLHxwSMcV2T1U3DwoW1PJOxYN5qBjwFf
AWj/KUiLLFKf0VMKF1BDyazFTOtIguuO/scLcsnX5U6mWuCYlQ/O/kwaeG/OZJAR
TCwBGxeZnScK/zCK7Kizx6FkbZLeM1yWksVOm1mFsddjJrvdJoReE7TXYaKRgMHk
f0y/vXRN40CyEyYvs0cOlgwY7pEjI7WI5nPASGgLakT7EjfSX+cHOYOnVoKMS70T
T25VCiZWbStsOb6soXkVs1SLQbKrzAkZtI6ElL9v6WLj/SAd0dy5srBI8soou9QQ
MRQRVYpXw+pa+bonux1OOKSTaFtXB42kr1bizj8HMYzRQk3mAzaD0AK4H0qxf8vV
Y7QS6F32Ij9lvEEFECzcUW8rc9XKDTTUsZdy1SDP8D49kzOYzgo7tIlFRioWCp9s
qbsbtpB5ZTeil1YL9PHRxvz6KIBTyEvQSQ7t9eG6MVw1kVtOBOtuRuLMrSbwbnFi
aR8q2MFD08aEB4c3cWkYONQC96OmGUa2tvRjTDmFFIBhPeofrGm1wUXTw7QEsesU
kGdbf4TSs7/Cqk/H84W85X4f/zBZz126yW0aqgMTWQK6crxWEG0hFe9x9EhnuXYQ
fS6t5Y+bkp0iVLaUvDYHsENJWemg+DgOOcPFhDrMP7AB8SeHTL9B3UFjIH0EqK57
HdXTd/mDd+aBVCPcn6WiFmtvYbLgWXGX2hfarUdTc2nkleB3yMQaJuB1JVvtq7UN
/aTYamDw5lXDq+UqrRhTucHNuI9MBcdYUe7b4n+RiO/mOZy0J1njSzKgi1NhVBAb
94L+nXBgaHWk8Nyc8aCJffJB/1HtHYX8dDhXcLfDubrPeu49omtuGkijuvwfH+nz
G8fD8zcZJnpUMNUfnwUjPu2iPxZ3eALETTp1WkUjhz8Q8LByjEC3isW0+lmDvSdW
crqOKpn2LbqIwWuutztXxyjxdSgEQJTwSkbs90EZvKNjEevbp8bt6rsR51r4MNZ2
yzD1ePaypQPYhyRRK2HF/B2X2y4kjsv7rCtDwOmgfecpdF6l+sS2wfOu0cFkO8wH
DppN7BRDmfbS8pEZbf9zIWz5RreUVK0IseHY8aq9Xmm93pg4ojeMCqbVUsvckanC
npeGYXgzK4qZcAfdfDiRWyCbGST6ibePoZ8FZ1boQhLM9queP+DVXoDaxZze6Pj8
aNib7Ac4gM/IP1WDryxSnIahu/i69dwcKQWBIPpED25BujrVHY+NljiclYKszx+Q
5KlXQjeI78rFrZXZiHYPS1ubQWavD+v8Eac+Cts3ev843tWLUeD/ImCeNyAyxTfW
mdZgBN6zXKaoyDwONgIrcGsV47nclaeAt1mvwH8M8i4IpAK2L7Q7mWpIBPujk7J9
KMgvhbhzpzYs/Ew8BCWdaeQWTvmdfwBnDL7DkLAMjkcN/cBhilEvWNnVOyasMG4k
uReiGzVtY78v99aUE42o3ii7w8M5obYvHYptze9XWM+g6V8j162ajE75alFHY8vL
jxVtl44rbd0QSTJyIVzsvCSJ+/ixoFut2fC/8ZFxCACezcz4Yrpsfs+mcuN/wirI
EWMLQpUtmn1DH/ijucKihWr0CmzHzfe4O9gzt0ryR4NflVtGfyRSGToy0L8eJ7/q
j/ZNqD8XZ8p7MX/ErR7Z3da/MAUb5uIo7oBP0UURxQkfpFi3nWGsdMPE+wlOSl/f
oJEVm8opwmN+r2CW1ZVoJKnGwFnaoa2tq7b55kmWDGASceGM2n8aql9iw/AnEQ5c
tDszKH4MkxjqN8rHurpHJiS4ecce4zKBtKP3JFD5w3F9QsdxBaijECLsEnMSIC77
1CKlY4ameeHq4c3LM6MHmxeUUisiD+YFxm18Y2wELExmb4NIISB+kI8bI+5VQYuH
IgMuBi94f2KaGPnMPT89gypzfQInUmCzanmLZZ8hWDuCUEG+vij4dHRAMeQxQRCH
WCJo6Q9AlrsoHhF+SqOFMN25aLtYL5vNBfEgVxGYZbosUw2JKlcBVNK7d5YxJKoH
YYB9ZrmrbbqDBDDsIaIsW27VfiNgliUvXDPxmjHMnpEz/feW0eihJMlc1ELWPJJt
9mPHbHcNEEOgu1rcGu6A7ctJzXdnrZrDnhYlCdMAVmPbLzE64w487uN3D93NKTaB
WNuGy9mTksAua+GTjLb6F0vWK2rumlCyObFsn5BFBm2p2Cu6DMcfJhpgGHpBB8qB
YYWWIvr/pLjZ9CVkPMbLfRVNJ6E/wrBVq8APIqTCm9mFZH7Kg0dncN1xTj32CFOo
Em9+c4c47MAvPqMiGgDH4kWofoweyHwyd1nED9o4kChSWPlsJa61zVf5sCmvN9V0
gDUWXMrlxjv4rcS/Q0sxb0UeP0qoas7OSOMkkjHYmD64kM8s7jjYd9ohtvgriNuG
GKJD5huujb/coL5JYbCQk4mlQQuLIMXndLdjNxOTt8WIpGQ0LPqctWdfGP686Vku
+KduOp5XtHx0rLWbs6mfPCSdQc14kkBCxBnOzAQHt6fEDc3X+Tjaps4X3+GGmLrO
8rXtRB5MU0ife93Mf9b6RolShgItbiwS+UXHDNRlO1+tSxn3mNdyo5Wch0XqSbDo
mXxxEu+DnAJpNRPwrlkfU3M3pBEKnrv4NFLOU3vrfze9+MXL+uPNekoXSTHdS8s/
vuF9Ed0izVYImgZ0LM5gkVF1e3pzvLswOGggTdPIjU05K8HpW3Hi0eZxuBGXFeBc
uwWP/gzcJwCNabsGsbC+pvZOqtnFwpRtTCBTBBLeF8VmPIFFwHsGZJHfkIyhEgwa
OWS5fKpuMvMNYwg5Hoy2XZ1gjSDJPn8IkPZ4Mkck+fAmMHfaYccnUsZKBtUX4Uxg
quapQ5IbQh5IhM+4YS/7i9HWATzJfmVWfA27Wxn+yORp2xHTUrPsoJ+n22oJFLaK
lcszCPxbPiwNJ4ZVpY+CdraRGYRtK/Hmxg+ytGQB+CI0ma2DAiDaN7KHPxY4/WYf
9AsiJMF/kEEqSdT8Tt6eOzhrvVfFK08ntxirCg5H3mKx3QH2syCsaEIUUvZkPhFn
/1pOVmXYJhFdlEM9hiZQ3UNTC1C2ct0cUilOsHdRGhobqJCK9YZ4QCxh98uhWkBe
KHqfrMP75jbewN4+pkOhP8qvtfEXX+/BlhAmo+QL671mCpT/JSKkbAyym7qzS4n6
JY2o4GqVJ6iRJPHvLmx1wfJDqK71YouJuqhTq44Z6Mkac6TDJbX0pDZlHOxyynJ1
K5zwFru5SJVQeUwj+7wLyXQ+ygvLg4jtuFHrKJAB0p33d2zaRRTBSGsXSTupxSJ0
3NMezzZ8Tbt5PSW7MotzomnMJ0QnQ2V2VvG3d/44KUyzVVA+/yK5VuV43U1nE0WN
6OVAOe0gsP0qRja+D9MdjHbBfuaxDPrxOXOC+G5OdbV/YqqTRD5Il4nRAH1S0PEi
bTZ/7+2EsyMLK7exL2K+94biAu0jigyWO82Ngtr3lzG0Tc1xBA6bzsNrctaChPZt
PkN2ABVvAhyO50xXGDNahDQHk3QxF65jes7vwqvLqhj+CniqV9dOB3vu/wH2/xet
jgkfUyb7oaTgRfAF65vHHc8BA3Vcs0KPbUCvAc2Ehy6nFdt45KlpZ1NQMAxpaJmE
eXIyJBIXFd0ZTrCf8BjbovNxK1etSAD94vzyBnvEgHJgJkrkHMmR71gUl7TUVfzL
TyWJqyTnQiI87c9NZnyxMKQfoGSwbrYoiCQrXyuy06QOjRTOdAWJDjqIcyWdHkUv
jRQz215UnaTIaHUAFpOjKCbzSpdLmPOuG7B3HrPYQqZKcwXmcQoxKWr/MuMHvU+Z
z21pW7fU3IYgc6MU9Lsjhz/ZHI+zYsZTKQidEe9y6eTyFDj7/99Xrt9y0HQzO+aJ
j0Agz7yeg0PxHeFQ3R/6r8c0Q+2qeRwOv7Cr/2PFzAg/2yhRWHZ6dqIZP1xQNN/V
poVxQlbcDkgnJAznbK/re3VWYan7JMtK0c465Rw5pySpySqcO9nztCeMtxFBA6OT
9nJPYKih+AiajZbNoaxoZHtb0s13nIOzjlKIGdd33UYax7k0Ub/rZ3apKwKKtqoD
W9Agy4uC99VwW6Z+vC7DWUmqmLBfNzIEpo3BZFVJSI9MmriLLrW64txzXiNkpQ5h
U7RhOMjD4fDmgbQZMqAG6dS6V7wHGbnfNTtb7Dq7DtYD437nBQOZhqhDN89GSTxQ
TEocl2wSHIjNJEJQKCYjuj/YU/f3ybAmMLodjIgwDbdwoXYLSBhH/j7WEOxSGAB9
KRZ3EUEbRAb4kFTOIt9h4suJyssbK8M5e3PEsJroaQafIKmaf4/ztovUVjcoMdI/
gSPuGh5kbAX1Z97IjtxbTYTYsokeCo7KOqtqnoxVI0Pj6lTfZjWYlHP/IkdNE/7M
bKIGIk6GUTRrKRq8JcEq+eu4HYigrGR5dIz7e9GEJaK6OVhjwx17qwRAXkK13rZR
NImJPaWYvVm7JVGAo/1c+oMfK5xegkqM8d7vw9siom/603wW4OwZw80aVsuSAlEB
lRVDLEWTe3dR0DCmrl+mfZFiV4hobm6hDzMWkSKImTCFxF27toZS44y/R1jiuXxq
Ns9qlZet2EW3wQTDi+fMnrzXU9h//cHizIJpFDpdTs/XT6+lSRPUQhOIG016vxEV
PZfDBV/6rwk32s7mwO92AW5iSglVwhPPzzzPuo/UFskTufZrrSZQwyQ/8Gy5yVIO
HhxkqRjN7AjLbNlO9GWMD6fVQ9riHynfssSR+lztw5U07mg6sz5/caIDsWZJqZ2M
TLCKGoW+GgyGYGtsnXrnLK3Bc0dw+OJLv/311BCocs0cUGgUJZdDXftalGPnLkpS
ZeBMV3lDjjahw7KYM3Px2drKK9oyJ4nrUinzrZMgjARqDK9WRDC5GtDtG5dCt5ei
ziBqt7mtAXA4V8iYNqO8rvJZgCejaS68U5ITyH6pTe5TuJUGpeK0mS4MOzIG9wbS
UTahUAVs59Afi+dnl3rXPHicaGn0MlxlbgMHbzSODtDroBcdjIVAIoFGgIqFDJzj
vhSf3JBBShciwB4GSEIBqhEB/hd/Ov+tXkej20X6JIRQHXZWYtH2YWXitHFhIShl
wKlem/rNz95iT/S3McE6u4P4MNKOUq+VXZrnFaNdPkP8IplOKX3lh1a8XqVSd9Fr
p//4I0R0XVzjJtOfvvVy55MR/SjgfdQOC1Nfu/nVQrOzn1wef/WnyGGmeAeoP5bt
MVDTUHzhQW4EvPPLP6lSF+EAnX6VyQeNg9ZmDHZzvOcrOl5bvZUbY4IABV8bmgPF
3D2yo10HOAVnmrAxAIG+Y3PDNTkSKQnfqlJDiOTsWreqJSb2h17KjM8JEzHw046q
JwQVWpukSp5OIqhjpvNwyWxhRT9j4mFbrY1orAHmakawHgb6BgTyCY1MJPN5y5md
fRTO6Qi23Q/1pQoQp7gtv0baChYuszpfMg+/ZY+IPx6nhiYmyHej5coRzJdVut6w
7CEQZTPbmCltJh+JAvgLLZhqWT5Xgq3CoufOYNednwkXqG9JA7IOda+kRZpRSyK5
TIiZz4HO1fsIH2f0RFmrfqVwHQR1IqlHGqbEQMO7/m239a39M5nPY8V5V7lXyxgn
1/z3vy7VG7v5tKodKwxcz+HYO9ZKhTY/x+CaBF+5WtswBZrXbc059ya3sYXv/908
CGIscAQpBawf1t4Lsk5xjTOlqv7YY1ARJp2YAP5VGogP+IGv2VmJDo9sfo7AVAgR
FL9to6gH1Kwi+bcv7wh1pL0veaysnCNKzn+GKUKNZVv6rYRitNNRdEQEj7jyioPP
b75zoL9qwrhDh8J3/Y05qfTExKbevLxu+m241SrfydcsRHCf1fj0PsV7GMf29g08
WzzaiNe1cku1RDGCuSEY7SadUlbfytj5wzPZ41OngtX4XcLHVS1wW9SC6Qv7945Z
MKVyCHLUA9ZLzMldqiC5tbptVly9MrQ80wOp1l7qWCdsiplBRfE4eK4RG8nZ/Lgw
OniUvrOAIVpQPUgqJ8n6cHj1mRQ6Dc2XSdDzaXV1DKKjy+5LBy5bpIxQzcFPf1i1
0HlEgdwn5iKVqW4GmWEOhnzeVQ/ZQ+Z3z/ax0TNMaEAUXCjJeA14GUkK3teE5vcJ
+4Od2JlIZFTn/Hbj/qCATTaM+yQZOlojKRHOF9V6lWEqqJxDr7qMk1kFa90lWCxF
w/O9sDBhB6aZFwmi78I700uVEUOfaemsoJQuj4ZoVpMnMc9MSFvceKmSJuUaq42e
OnoG3/DkpKHHM8hx8wL6IZAfZn5I2tXmJQRmGlZGET/WpKTnPwXINh0rpNZXyZ+3
dX1jIx7ir5bQI7XnLTSwg5ICx9iNVlJhhipyWicdLAwJ4G1qPP1C4uQ7QsQvWTFK
xyP3xFwLRLd81tPnTvg61Wl4ZzZKfTIkMf7YM+0+ny24NGqEwYNPupZbpYqCAYC8
AwLMUhJJV8bl03w1cOUiqlDbe3PrfUC/c4CG55M7nhdMwO2GtON77pAeMS7e9chF
5DIrGfPGrlefwohs6ZOHNRC0TNsJDzmasSB3Wy7oqC2ZmuSXmrUjcKVlfOX1vnTW
/ULoZQqWCwi1iPRxmlWSMeqex9ML1qLNQIGMjF5+pSWCzSS/XTzwXffitWsLAiGQ
lRryPGI+Qo9/Qzvq+O1QgQGnnPR+fQ/8j3mtIb1AZ/HefQL/zPWU0XGOKIavzX4x
djWt8CXwieUlw3d7X5DOufU4PJ/ZYf3Y7q6MwqScwlGYZDNDgxCcBFBQ1bxjAx/E
1lru0xBkuNPVclS/pL8U4f+VASbm2okBzjUaA3S5+mCpq5Kf1UT621PbBZGSAc1k
0f6lOiL3TqqYJXbIo+lv/GFu/qUALqj9NXzhEk0vpXqH6awf6ZelKCWOxkcrXgeR
LSYLs66KRVjFtAiLVewE4EiYfC+lSLtLR/bvpnADBOEXa1qLqHE2/oXlCAV7KGil
z1Ch/iyfSD0MuzsRMEAyuDhRmWrWB1TPSBFZoJz9gjbcLqhTtk5E7x8htx/AAXdz
/+K2mKUKez0SY1z/2tU4NrjiDlQKV98rwP+pKlqAxwen9vfTqGqu/dqLW4IZurjh
UrQomo0b5mOGcwmhIZM1oB/hVl4ioy+TwkeeGMBqaccqT+lAKIEzsF06956T57Mg
/nJUSwRoH6brvHbBnX666l1FE8XyE8WcEIhCuUehnErSRvs+d44xIKBiz4xUKdAp
iNXE3uFiVnaeqZX2cg2KXampcqeAU0wCFC9wheMtm5oUkdHT7q85OH0gp13aQeoM
ZaWyWkHfRg4+dwn1hHUofMgo6VcLYCEu/G622Bgk1DRAICi38+BQHAbpTU8yJI2B
N8E2iqaOSmRVNWuApRdUDPNow2Z5dtX02uR0+TjwWMUoTnYuRZ1WGiCzyH30F3Ce
YsgXqgHeA3UHbgLQ7VA0r5Ax/RmPJ1Jni8/V9gP5nThRh5QTomKjER2mDA2cdGuF
cu3U3uTpJ7BICqjh6NGVmOvJWxdN4aRDSRKa7njV8AtT70oSHq+eRFfC7Q0WTVlZ
Jyhj/WnldYm+D0XEqKzMDbMngPmtACVLbbaJ6TddTlfafbMma6zMTpBg+NJuVFIp
Qd/6ZK9qztc63K0t7syjbDWt+isj5jqUBdk31a+o4AfTNDmNZws4vzblLAH+LXc4
bohhnsasZJHUnxeGrRk1oJVtq/af3we2DbmQh2utTP93EXZOeWIE8sHiyoN4mAtP
UmT5KSuKbPyTDbRh+dkhERHlQhxqCCP0lBMAVHfBJ3/jRZMfZF63DD6p/Ca7qu1C
or8XLCDKhhjig2KjzEx1fkLnq/aHExMuLGiodB9hl3xAFrRfcV7PaSa0l5zx+Al5
8q4E8v2bPbaaoYLR9dOSL69cWH4rSVDDMgzyplwU+7xbl3UIPzNUq5Pinbm/kHIW
/mGO1BtjFwOc2yygPtUYuD+9zzR9Cg46BG8QuUEyPW8FqRZfnWnV+PXIty9gl7T0
XikLrGpJQgfvQAMx0hDYyxiM2Il3ZVZCtZCAdgmDbiIxmcbMvgUP0c5bB78MRNuN
8X3zxDwgAKwj5jwXhcLoooCnD4uzu/lG97Jw62kSkpRjf3UyqJjwvnaG9zXqZPiN
twj0atX/BsIIm012cjExov8Cm/v0OOJASGeYdYYJT0M58PQlfQfD6J/E1IcftXg9
IcQ/xhHaiVrMYcKpmfTfUEIDhZTWHJOcpdM/assHlrI/E8MiGB4K3ECRVvtOocbk
qgrtNQN+zX8B80alLt4J5ocXeSRh3v2tnFricoA1Zx3ZtG0ykYGirrxUsXytbI1P
l8cwoZNTyomMiKQOhfd5Q0xsX4rH5E06uzGq2X4+CXPuqDmx69pO8wKBprzgBDxe
J7R/ilp8aqVwMBRhPujgLvpEQe6g6+OgmFitwyZiy/n+vTkTamPjzpi7wjLFEzpj
AG1ZTiAwBe/stnLzjYwettvjHXxLKxqFj1XFVsWxju3o0Te+k4o+ZHx2KNGYF7Kf
n7hXntcgN4Brw4Dn5m2zykWC0lS9cHzxUwkDN31Rmsspp0d0LZr+c1I1Oe6QzF7k
d+BRasm4fW1kd6sLJBlcSggNxheM/NnoKVDCVNKDr0dcUAnHgCgragb/DgMv87MN
DtHjafrzzXq6cKCOEJvLOQDWiTOF8+Ix3J+vXTj+4qAOQ03nQ0WhI54YMbgj7bsZ
1vZbECFiKatC3CeSJp1YRVPGYIt+lpH7EANW1GRbwb8RyryeJ++UosJ97Lngb8Jw
ERs0oIipPG750sCLsCX15lGVYCcbY2R0V8jrIlHzTSp1I1q8QFPW7tC1jigtlVa4
zFTE3CsIf+CU+x2VZ7gGX5IcGQvRyCzuKnvP0/Kdy+W8c+Ti/UC1T/GG/GY98Tv2
izj0Ee3NKibXB5vvZSu7/PsA0OvSleOys/GDa6LunKFgNCe2wHj1LM5n7M/4kfMy
KrhJjEJ5GQ8erGTBwYJzEUwL8pq31rpthBjy6yk8lrRhMFKv26d829HDkcQ90VzU
O5T1i4osgczdQ2v6jMalWnk6rSqgNJkNNA4JIlAVGjrEPQ1jlGxZMr1LwnXr2xzp
RwFG1iTiu7t6o+JdUow25arJ8gzGm2nZkpqSf6YYEh3hKXJiVBqReGgPmi6e5TmN
AqHRrqukFiztvjFBhCF+qGrB22Gyz+V3qS3YOqcF+bsSUEFhUtDwAyTdk1YdYmN/
aeOeH5t0EtbFauv2HyX6iix7pCjGkYxF0kY0cj/MO+nmRUuZUVO5YTg0wYfeeXlU
30QUXc5xwWgfbbDXC5EtgFX8ubRM++6sunqHtIb1W5Y7cjg5nFWopYPMXr0M+14f
lDfXZv+oeY+Isf4e8vKgTA++vpF16fa1zLmkKtPd72ZLF3defoOyGbs73YYsvLBM
Raip4TQnANylC/acTD8rxlrLkxXfJJQsn/YHEzFhKb23MzMN4nTEjSIIZM+aOU7l
C80t6ocud9crw381RrFp+PO0VfPTVSjdQo1zCIZdu7cjhj6cAtmoouiwpJLhDAPO
Lhojab5z12Bos3Inz3EVpKpbLmI/FIwK1Zpm68vMyTMMWtrpTzcAJLQCGSVSVY/h
Vgy/y833hu6NLuUXdg+eN2g2BWqscstxoczUvvX0DVoX2pZC9kUq+8YbK1YYmYGs
kwqEokHZxrm14GLLT+ix7HqrGSOngelxuy+MZ6fsQEcUVeRFGhXBqzlZLLMdL2Oe
JDXpCusMdrCbNE1lFDko6tN4976gV4I760D6VaC8/as6MGxA3ggLYBD0TDIGMD1X
wtUNR/jH6JNyhns831Dj+XuC03rF+NRxzxED6Zzl4dkQlYlFRq6jES6unWNXc8/N
dFzPd2iDl3cbPK5cJio9WBi2PaZQhp2nAZfEsT5oYdnG34QuUfn91RuLJkDEdYZ5
7MxMZPHh9gWXv0ktDPxfk74KFKqA2sz1RiZb4Cr+qc06XeDXQwQSoXVqA0KEAis1
H8XLHsEsbGmZ+alNrjcaHku8KAMNISJlY5enUAY1/VgiJ8PuOOKXvLwXFqO3bQ5u
r7d1sMCmYmOoIUz6daoe42lKihACWXcj4Hc9mMaLVThy62Ti0wZfzmJd4K1AxVPj
9eo+wEu/BHGSZAV6jE9ouZuYmXOoKbT3RTNE5djzWergYHkmU+pg5okCWEcwLyfD
zJHUsSULxTMiEFgt6B2QjzC/Ff8qDdTi1wFNFxYir9Dya7KOvbcc5f8eoJV4bwim
jN3pv01Bp7+iwp/7hOD7MEQV1YE5GNNLhICrMtQtQun+E9MG17/JFi0yt7Yra8oi
jEE8iFffy2uTH9SGZoVNxIV8O8Udc0tnvZM6iu1nU4MbPNBWGtzKQyVnIbj2LVxv
wzdFyYbOGpXVdlP1OkcxhyI1QYO2+XcwFHKt+WkNXCoKluXJsUWW5yyGacLcCt6C
amlFTUZ+z/M0S/1+mDDOlDX03Hpo5ZM55S8bXbo2I/sJ3pku+poO1xrwQ/zR1A10
aFvqbqbSphIrZrzYMf0Az1mRItI3peMYt/pavUdqMdXq5j5BfIKP0Z5oW+L4kbJy
Kr+Sb/AF6XaveZixvM/66O1Za+IsHUh5zokv6CyT/spaNF6tVIaF3Fv3BXGoS0TL
8xSsxipLdXWHV0h8JGP10UaMA6V6qSuNkaVEmzKld2cEMQEb5WHOpXvRf/ibscWF
EJChXpMpGbpnRNnEHWBAJHVuIyUmp9wFiOb/iQX2JAz9rendtc7Btcv8ZtoTFF/q
N/FU4HrAfJWoVHC4/HpE9N8K0PIHGFC54eGSs6fisIC7ZbLftUyYj8S4us0ZMP0G
/0laf/ZJlY5VhX+B4Te5T90blt4jdAfGIKAddx6aAb+eZbK240Nzog4IC31akrbp
bese64lzh7ekotzoA6+sXywcd/sNxWTOff7PokPA4LTdbT//5lG/oBvo0qtV/opj
aLrYZqcYfidF9xpZpMM+pf4BfxUe+BmvWn9togWl2e5Bdqo+p891ukJ4Kc+NHD3n
comKGwakwhpujF7CgNJBboVdI1U8ZvC+1Vz8qpMAaAzkiZBPaWimznC4leKgZZPS
ZfrpPcoNzR0FLaVPr/Aa1zP4Ygf/LEdXH+JjFpYV1AjsZje5cdfnGLCvjtCSAk0a
pIVSvSTuTLl5DKUVM2/6FZRyXLQEQWJ053gOPePhDfQ8hehMeNs1wKzgWbqyI7VT
Dn1YKOnH6rv3dPemmA+CKm3DDJ9bSHo+prR6QS0gxo+mTHQW5/XfSSVVchMEgk6b
yX2YWh3xaRwxKZ2ZtVfHpcT5Q+V1VXU4FsNai31RejghyzQZwui/22p/KkxgLpKa
tXoNxEPFBE52jBSjRKU7e4k3pc+bwL6jF+Dc6P33YUcrKFFHWJx8emFOMyTl2OYe
2bu/+MH/fXPgN74SH6h2Tw5c7tyMSY8TietBZg5QgMRS1gHPGHwd8pa2zjgyEDlU
+DrZQf6JvI7+m4Ct5NawEG0BeyJkItQO+gjhrQO2YED6sZaSiJ43w3vNSA+JdPzH
Hz8z9pyDeWnyawdhT343v9ABpCcUKKRijHaKDZivDqi98ibA8RK0IGbjBNE1bod4
asOYDw1tPrZTnronHO+kPH+IFuZc1P1YavlGrx02rY/V94D5+IvTzMgQ8xqvDX8I
fu7peD7rH4Gghso2P+ma3fAV7I64uOGpF8tVVYsBRPnd6J6vDr24XmPlUG96vVn+
xyElkrrJMMTzKY/U1rJtSVb/Pm4h0X/5oIrBXTgrjIrPYACLs08MoexdQuZO8Agz
H0+lkfenpKDBjpVKp9s74CpsMBEehZ9z7AZSxGOioa8NWuxXhxl1+aBcIK65H3mJ
ZYNrMf8uLD248VJReOmTT63eZOC8FfIAm+cMOQlKpTNQiYpHVWAczFNeF1ldFg+y
//k+Mk/ceSetePVvH59E4kkv3dGSPPyCIDQF25Jkzu+bNREoukPgLGMVEPjJw4iv
jRGVmKY5zq/hjrKk9+Qv/ULjSqzSVXULojn+BAh4dl+WJ6FpOonx2OO+Pq/6l8Gy
Sint6CXpC0d46qX2KL/H9st7uJvkTt99RR5lb3u4Cq85PZY+LDNnLoYLDRheMAp3
vv91KRyX7Enx/ObvbVVxlygsmjeA8u1UVC456BJJMwuwQrbp1CXwr05wfprGw2rx
VhnGaFZzwb8tskgZSPZ3vmBGBUa8nozkSEMoKpX4dfiv/IjErEjxPgMOsi28rfqW
+veMmE0M2eUaIVZpCaySRpunYk+/5Ef6EE6IkvvvNHySDner6nO3gazi2vURe1Jy
eXW4VwKSyvcZkkYq/wwvRgoBUY+wZlRQpN962Zo7gaEJ1QYOjlevHH9/jwFntqh/
6WP8HoT50/+Vkxrd3AUJlVxCSfQbQYuvNeUjF8G2IY1OJlLKoRU4Anov77e1JHtd
LvwBbPF6GBowzSF0DIm+uDa2DsmUmam++qW4sxOeUELYdHPzIo67jH+ZUoCNxjSS
JleDiRhv6rfpXSTF9IPSvgVQEsSzoHznCJAlE2zp71zu+4ZseQzqBSqV80APKgnj
0YKYu4eEImkM414Z/ceScF9CLFnxEdlHWqwoyChHUTTsDzztUsQxG8kgP0SCRLl8
tD5it6enmSTFUEYIzEeoOrakzCqfOcOtrOSo1ed4P7IsBtYdwhk34gFjPZo/cL6I
a1BTm0ecvl2QYyBt7aGEYWTnlVsaRnUEqj38JE360vNzgMKeU1sndLGCTrCU+xP+
4AkAHZSc/s4djNXpHetAat/Cqy8qNGcG77fSnJ7BC/h4wgCIjvsIvdbksNhfH4qe
Yqk3uOOEHxpJypnAtj9sWsvVIzkrJbxXKxsYeyY8wyytHnzKCbdDmsKkwdiGI14Z
AzJfEaDQVI6+kGrAEcdQWTgR4tR5gJTKF2yv9pwssmHuXf0EPfrpkB+VUD+9y27j
IZmOhNtp3WV4QSDITQFW5BWBhUNwcgNZHLGT2ZB24qoRDZ6XD0gf689Ve53Op9by
F2m3vKfhn9XHOOv87oiOgp2RMa0MXVrFvlNPX65K5PeHoCV1nYrtpvLrRZhkyHH2
nWDqRH1aPWK3rUhR/Cdh7RRwzQNCBqntbDbb8t44olNrDcRwV4pxrM+MyVUEN6Jc
DEpz1xum/n/dTlH/wZHNYk+QyQIkFT90iw9DI4KK52+xSugrZteBnTQte2BJ8N93
BKTERK1fwC6+Ix6nAf0FFjkDdOjFv0DWnHgAsJBhPrt+Mr58rLQPMrJwU2lo5WfR
Jg6sYNzhV8LYnlX0gLsbgTLGTONgRho2L9grSKv4Ge1Y+/gKmxGs/r5geAOpyp23
4k8lucEFpqwVZS3psBrc2SAae/PCJrzntAWWlioKRxPxaLeNsius/43/X2YNxuCo
iUSiWn6ad87L+g3GiP9l9/DHHsxfydgyoIniEyo19XgkMcGTe93HHKr+UvxjXMmG
Vclq7pFt1BzepOLNZ5mbnNWiAKKZi9C5W5QeZlKMLj+wisiE41lA6W4Yznhi3MYY
bh502Y2J7kQS2V9xH44yhqbEV/yhBssTdwMya12L+9ZsplpW9mc+OIMFdeFrxz7I
cl+LE0X7gNjczOHUnwaHPENGbU/Nnkm6SjTv7MxfkSnAR2Nitk6WOj4Vlj8SVMXJ
pzP2MLL+SmaGntaISRqS4mDNkm/tHN3IwOTuZXS6KjnmaFTsmSZxrQ138oPTjP9m
9cGUs5XLWjaaTMzW9YOrePHCtRfuUUJ4hGuoP+Ay8p4nsdf1yz06su9uFBb65XeO
rO5O+1LqKYFnstZ9kC/hFLFAReWaFNhcdmG9lm7YZOUh04TyJBsd/mwS0TkO9IeM
b2lOS4TvzdcGYVgYHlWTXkY5N8zLp0Sky7eA5ZsNXzTAWC5hR4VGYo8oXgUTYJwG
OeDR7t6mAARuQQPIgeHQZ3BdiPFQ6bvQhOM71mUrv2C8sksnyAF6++ntSkSGhngM
gMvUoK5VHZM71H8433pqpeJo7f9EPqBwlRweBdhLQDvOn49EA0naFoF3aeW6OpJt
h3bfQVCQ8lMUoFxcMgUhdFj9i5UzmXFd/eK+QFUkTM1a+TiqYxFAnkihxaHtg41N
nyZz965uoVEIfk4lKpGKQIXTjiR5XdaSOfOzX74VOKPp7bYOCQtpKCtiIKDl1/Lv
mpkiKZSj72wk/6fEb51+GKgrjdugwFUqNLBgmQsCHHEX+YJTCqnoPLwOO3jSVWbF
0lJ2ohNHp00oeUd767c6Dq0/8d5s8rIyFq1GaYxtkJ5CteRrI/ScFxJojMzF7daV
R426PYmYTnaohHz1QVZrBL+d7PQ7jHnlu/kkb1f9eR4tJYEAJ9Hfk2JG8hSGeFRi
0lyZR32vEwHfGOXE/oW31PTY6TdXDq3oLEDEwZAqk7MFx6qq17HzSziuJJliG/iu
NApovCnfrW7UT4hXtVhtMyOzzALKWf6PhPnn/4R5VbrM+JyOiCld4W4BbJDC0UE9
gdzKAvtDPt6AmExOrJrREz4JbBKctEGSJcYCrpfcbQif/MFQl0wbKDAiHez+T1EU
G2Q1YVJD7LAVV91CXIXEBkwDlmSuVohD/yiKBNpX3YkEdfr8WVdiffJo8gZQ7k7b
sZQJax1bO3HY5SvN+ZwMdBp3BMllGpNVs8Ewh36nKuq1q8qvREfiiy6ZMph2p9Pi
vO5+81ux+KDv4VWHMAi8HMjpyKjRDmOrHrEuFFE+Flp+1K5f4mKY2gVPdrIV5ZDb
2BLiuHlH5BPf9BLGwGZZpIKvQ3iheO1PzO+QKIfXTkXFquHFs8DXPtpwrOMD7YIZ
julwWStPxyiVjlHP7PFb7IKc67hydyI20/dEk55ZvAGr5yDwq58ST138Lm5DInwU
V9VVwWNPpOziKx7rCFt+Dsg7de++wXMUWTRtsuVMNXmAjINa4sIIF335C4xmMeYH
NV8TXox3MwiuXSdkRon8U1kxVGHE9t7Em37Hmxspmq2U/JasgXbu9KJjO1kILUee
g69ndM7nczsNIAvLNwKRRmTcjwz7nhx4TnHyRRWpNanf3PYR2KVJulZCX6JFJcft
kNMjft7zRgwlPUu2V0r2krVTPaz8oFarlEQ/WE/cRUXpmAX5d/5cEVPzFFcLWSKr
UBOJYgWEUQgt6kTOJW5CUfTbJZ0TKWg/UIVzTWEVckKo5YPpVhidn+xegF3fvs7v
2cqOT+baC3ufXw7N+a3T/juVlBvCsB9gU6dsV0I+JQ+5k664KtteQRgkAFct0ZPB
/6L0v26SdbJr2aJWnovvYBdSB3IwR/fbNbSGjkjnlA6cYsNUpkA5VwxRcXezmq8h
s0UGF+bf7KKhQ7wlLOI1T0K53uEk6TEadEey4baorUKSZ7mNs6jJX9ZxeYeuUoYU
/2nT1tLmi5CJMRXZuzM7CBcDKeZvEtcrFuuUin6+TLeDKqmrnZeeUAbWHGikHxyo
WJnWSS4Pc7egwJDeifP9B8mP85HhSvssAi7HZzqm7XpG6iQV3+PgA1Uxrm/Au8QZ
r0rep3xXiJeyTCBAbZFu2L3+RG5YxGPIG6nDP/iypWDnSdiPHDbDMKxH0va+r9iy
SSKu1pmRCZ98tOv2NgHz2mJHDpvNwqdhVNwff37/P0D2CC8Jr/aGwFAoPQn6Ag08
twbcUzMRFTSDlM4qq95ptQN1gPFQZKAfmT0Seih1KhQfdG1habTHDPOqJGuSP1X1
3fnyIdrSXWjXaPiwm+5JoBh2Qti6yoQMtT3K5ZhWMNQ8BdSCibPx45CTAFlLHQiZ
DlRiZa63YpgoKOzOOscCZgWjwUIcGU+fYJy5GksshoDC4AUrKUTp0AXfDWWzHv2Y
pA05vK/rSxFgC5Yx/8m0UEO5SnQUNM0yJdbd5pSxSLIR6ngvK/V0XMcmbvIm/j+H
Db4FgzeAVUR9n9gzhiCRFrzk6/kBPQVY3gmfdRXm574fBHorivy3HvCTkvrG7yrg
FBL7SXG/gNRXP8SynLEjj8T7RWtUjTDYnq7pfhZdTdeZf8OyKNwsw0A+/5Kx5VXA
lAM6KeMZEz/6fpaXYk9IZngub3u/Pwmra0kWCBw08VduS0r3qTHbegHADiy+9Vv0
Abbi+v9/8aypNwgRgpCnOxgHHUTCV/EMOAWqO5O+XynPmxztH+/YxgchklYBqBbd
c17/l8X+XSjbPJ8fv6rexVbVlqzharpFdTnMz7t/Sc70o942ADmX62jJXD4Fen9D
KOcigOm6RATPUfhRIhXEc0xZQJCgH8YyeGoomXpoL5uv6rk5neSBNSSj2FDqkBpe
QakqNH1AEkxIroyr/7DAV3PLDctvRZSdMxRifMfedjZAl7Mkz1ZFHYLKXg7xd5Lz
elPy+ohOulKiI9iGwdjXcXhbd1U17xlrrRR2eU1wX4de3tbgDzxbzM/2Sc8gITeI
f69ILc9u6J0XaBWX2Hs+IzY31G7zG6IOvCp7+yiOAto4vsaYGDEn9iWdQAD3V/7q
iwrw0z/Uwp+ugVs+M42B19Mdj5xhPS6hgjZAW6W1+2EJaiqKtHBWrSoEoBN1GFb+
roKWJ4BdfxT3LjYtUYnQXPkU0QMJux+gyU5GH+cDkbu06JwO0IMi1IYnPClIWUaV
tee6++ye7DfliS3eFm5bTCwMaB/lICHBa7g9VvQkYC3EJFJvPphAONCCFb5Bty5O
TEukhqSd7SIxFIT7KBEVykgavYFcDNWVS0+NM6FvaH6reOYVnBYv/7hetym0SP/b
1KW16Ngik+5tX9m3iXOe+iYyX+LWHzW2uPJ8/9xRZfIatMQXcpHpHzv8SvvRHt9X
nlDmd3MUQb90xzzUWwJTAF113n/9A6jndBxxyxBQCwcJ7UZLmjnMV6XHK74km85J
yB/Bcys732u5Fu9rUxYtiiByv9DmFbGHlaFwU5Cp0fe4PhGZgxny33IeWE8xL6NT
xOhXFmy1Z/DpW/+m0DmiaS9yBGksq1Sox5+V20iAqsaxXc+g4lIj7BOomEas/7OG
0yMk6RuDIGjcyJBhXdkC3kkywJsfgQ0n9+EZY5grmPL6zxXZ6+JczefDuS27tG2u
UfzX3NoddOKHdwFf3HwgI9tCrjLab3LMggrPc2VtYHYFEDELtTMSjZzcXdYy9JBj
J5/iY8uaVXS0cxoyrw9sGVST+F+L89Lj/FXYLSl0V6+ZBHVFnmWPSZyCQuuvfasb
4W2CnasMqjf7Aa3wEAMR/9+vMeXnSmW4kUf7fiUhAimpUHMv7XzhJA9Wzir50LtU
VD7+5iNQ+YucgKnUVzKduF2vMbH/4DRAk/A1Q/AlY7vkRkEYUg/q2X/4Pudv2Q58
f8eFsUXUKmxRJefWBVxSM+0SOvmCG1wnE0KkZh30XkNXoUa0O6wKa3DUKZOQ/fLM
RhblrblLazPOmzmVQAcdT/I/6hYqZ5tJprAO6r5I4pdF2u2YIapz8Q8+LTVd3XxQ
DIXlfCTH8h2nm2xM2W5p+91qHeHQby8kr3XIDaq1sZ+K8E4+hVEedt/3bqXtWv7W
3qxb9EjW0L+2ytEcJmNcLIdkI+oWhkp1GDwnMqX7AYnv/s7iq5rGLKK+HYw96zdM
rQvo3N4smS+0wItd/fePk7CnNO8B+7VoZyGUjnwchlyJpep029swTjO8pXtL0Kvv
jegGSgZuFI+9J9vEh6EmjISLBELSfB0w7HmioviLD3ojh421ULxTeljTJOmk3Ucv
oQqFQn2JZ8Jzq5Aas1mA/nYl1/x0ootRl2DafqSO7YpXz8OVVDX7gBZJ95Cs3LMC
C1xHl79ljj0hN8pJRnAKeRp/wUeH/7eh/nhVcyCkEd/N8v4JWVwlc3tIkPMFWrNY
ZlQhZf8GfhPP78Mknje4aEwecs28zrFKg1Bpu0ZXAxtWIK4BGXtDAk/sVPlI4YcA
ClMKEpvG7JsoIKv8Tk7rZW7XgGE9DTgjGPZp0yFbsl2z/ApwGEBZUUqA+KpDZFmz
1tBiMPSrujLf0FmYBqBnp17Drl3vCGL6jI334QNu9BzUCgqeidc7z6jTaVlyKh7c
ApkzPRZlY/hwr0WdJgODWNF2bZzN5jp3AADlIURdQjNrlfM6a7rwG6ifPmM7AQc4
SzOOSxQojErIwZ6VY/AQ3AuuCNp/pA1GmXwraL5yH5I2O0KjBuMgGmZg7AxsFghc
ehik9LiMd5fHeIgJrcAH+fzFN95DXyGoWO68CmiJ/DZcpVJd2aGuJQO+P5nfW2Fj
3whGmgGHS12FuiJIBZUZYRc8ucwMl2dLc9GrwhYEiIDKFgkpQXfoOCLsbo1AfhIZ
kk/a2126zC2YSGZ+zLKYgIniT3r1Q94FOeYV6hjo89wvqvh8tmv89iwHvmga50W2
7A5d/qhFjYbCQjbCFYw+prjcmaG+1NcJbH/k03sxIteMe8fkrig/1lGldgW1Xk1e
TQEU9GIaH96aqOvSYvnUyN3O1MdRRAAgsFS+mFl3pugLesJFePVn059HTF4WLEeo
+U5SOsy3CSI3h38x3zUKWltzf9JbG4shG1UO7W3kuB01p7I8U0ztdTXlfqfGu7va
vn+CiR/6ErD06F/StEeB0sgiHaeSOcX+Aht2zJb4icQFGD55RspgtbC9fKNYur+4
nKPuxEv0c45+arDOpmwwMb3p6VQwAOVCKGHn9EIv48GE8Cs3xu4Zxz5cUUT9q1Sf
nX2hUndiJuIhN2jqJUFFsjB+JSD51JM8gGMfv1hGZuPPfW1pO2n9sEUVOwoWOw+b
aw4p+InuHjAYQxPdhcets10qCvQbXvaH5rSJLqYdJhMCGwp0AbFShm9QU5yqc4vv
R3/KHOXbx1Y5QfsEt2OW51JNBap44FnFLsdMmnzusYJNPoQhX3OdzdFyZEdOJGbO
dgnwvpQbPvf9uGb4q9uyP6RAnvnOji6PQ2P12QN0XFNY5yhrFNnGqhWZkJ6MyHgF
6QosKnN42NzfLzpxtVu2SsE4q8DJP8rekYasTu/STan5ELQqQpgM4JNQ/A7IWHBa
W6gDLQjDJvfHVzppC2X8C7v/Jjh/zCebTox8maVKARhz+7na3F1mTLS9fZlsIY4W
kmOPqAK09sPm8S2iN+l9pV3inNP3DsuSBKXcmZ3wRmGK/Q9OoOPesCaN/J3Q4JSe
PlXLYgVmIGR+OtC62cBeOwh/5zRA3cD2wvrWJSpRY9hujgdI1Za2Y7siWINl2bmh
wRfarXiFs3NMFW6zChiiquWpg7NyZRX1jIhYsbjHa9d+6l+CEZsd8ka+WxurzIQx
ekUyF3QWlH+4AEyZSpZ3l3/ceEPt+7sqF7si80exa60+U6I6t2fEa0FDr6ljvx5h
5qiEiVh32zg0rH/MSazp8OzaIYeqUx0FSqp0QmVml4/f02eBRqZpLm+gG8KfbUIa
TEGkvI6a7414/IaITtz/66jplT1kTIkL7F3e/mth7Do13sYLv2wkFVmAqMfLErVO
2HTPUn9aC+PfSGvZqUKDzVTu/Yfef9XKbtaSzjdfMiALYxXt3XPElK1FuhawLupo
JzirhKVwKmHtsReCq6JMQ3u+1MBHG0UK35U/u4p53C5WrRwJOjvPYVVbl7VZUHXv
xrOvtSQpDLrnzIvCuif8KAcDzCDAkjRxnsI+unFTxjp/5ijqtaWKrQYFP6MWTa5w
v9ziOzyvxYvG09CPUG+4M3H2fpYVix5f/WBi2VBySj9MaY1W9BnU/I2L3mKLddSE
p5HlFmxr9LEl+HlfN2CAnikRJdmH7+XpDJlmj5rJ3xCxIwiqz1/C5oQjEdo2jDgQ
b56lG7OlVPqDY0Q2kn4S21UiKXGCbNXitIPC0Wx0Ji+8PTAJ6eu5vAVH3DnuVDCn
U/sXuni5uTUQbi5BUp8IeJ19jmZgsbyXUKz3aTBep7bxVG/JgG7p4K3ESljWzF6j
vMzi9mrmCQ2kXentZ6H5Hy2HE72Cr7P67fmJv3abzFV03lu4cUPr1F9VjbaIsHcm
VDKk9scTuLQfXhODqFg3aDPI55+mkrKlHGgFY4kTKkTjCbPWsV6ugMrxOEvbR0SO
i0d6CHZc/T8q9hl3RvBmOWC5RsOBp3Icebki1Xr8XXzW6Yvjm0HjMpwCR0J03JXj
JCIenojbYlKodus8zyhHJ7wSXqysUGhDwKTgpCQTHCq4TrTlfV618v3dqVOuPuw+
fx7W5VsMKVOvgv3oeldxu/131+8ve+zY7YWIPIJM+jccEu2S4fxRumX+jYx7LdKL
ec2i2kESAlPydqu4yaNPpuu6A00qjyH9yfbdOqEp3VIlu6OSnTOxUdDG2xNeUpcd
d2zx7pWifNcjUnRVlYZUsC+qGTcdvmmZdr4zR+MkEu6P2FVrjX36bGmHRaTI1BiR
A+LTpomKHGEjLqkJYDw1+/PwjhF4x5EskcgvVmuae0vVqkBzWa941vf1flerxaje
9VdWixYMKpfw2P7KZdLNepmvnllYOngjsiOR2Ls6EoSAsTKAnh37qhdR/quBT+xW
0oFrw7TGxbEs5TgV8DTEyDUUX3+TpJGEyXku5apg1+rg7BJ6FJs8LKAFAcfRKCaf
PwSCzC6qCW4+a3Qsv8YMRZ9348dS1o2M1BjgbDHSUo7kBb5A2dGBOHoxtFs7M1IW
dtT90AVIS/IQ4E4j0A0zTMWtRbIZREmy4Kj+6xrjslwCI2bc+n30E6M978wfmyYz
rifRHMlDXdc3cyUukEeOvJ4oJQjLrRybM9R2HvZZOySqZ44VNUjkIZyehym1cyJO
u6MHLt02rqwTrKbSuwyvmIWrjKSSjvfEbG9/9mTvTA+DkQexcb1xZ1FdX4/6750V
bMCNFXXUrBV50fut3D/xU3FBo9kK4PzL1QqdXSTx7cz3DC7zEr/a7pe7gCqdBpzr
NPktNI2R4y6WqHfPD8dMpdr0GD6VGEPWzQwV2lPXQ7PeJs7Fd4szq9Cs6Vn/AKwE
65sJp+IDPdLmmU3PALVAplo39Tjwx5pdC36Stna3rgicmGzitNfI/L0nJALPIDI9
bA2PZH+03aHs65vhY0DzOHLqp/O74K4iT9BEslmqstx49Nk5tCDyS2wT1tOOOKZR
koxtCoSsrntzjv9yfmPhKazbUwerey0CCdqTLvfMNb6AF4N2y/KkzmR3yvyTLaSV
pJ6mFDQx0uWmRMN5l88EOfttUbSUrmggjEnRf+/M2ik/qUZ+hMmiR13fPV1Nbxki
zEHPxWNLgOSBO1auZc2xChxPMk3Uwd05QxNFeLPpuIi+5ENrsWIOqi/Z+FwjM2lD
I86e22kK6ZAE5Z9tgTx7CSv0l5yNXajBJfRbQhdWv/dpmNfqUhzOsxcebD4qQKRV
dL1ktuOUmU3gdmdWUBHLYezXYb9gUub8+sQDT086TVfl7nS3v+c5cTVP5twtTOJO
kDv6XRNdIYdwW1hsyapJ0EY7mWmo8bGkN0HH1mPQAolrfk86qqdkmMoOZ+7d3JEn
OnlsT4qJV6WWYgAFc44nNvlR7Kv86i5Z+VJecm3fYDkfu0frm3S8KJl8R40/saO5
Ya25ZGYuLznqTjCiGQvpOv0T0wzDS0NKwno5wbKwjqIiRRw3Jr5gYEggmBtG3jo8
lDrA6abhBu2j9SQN2TO4NQFs7wXDfwVAn5mhEvvTKemy5IdJJ7ECMInx6pinWYKb
mVzSYSFlBOsupduc4vU+lyfloKBnms2KKrA3BfUxd9fTZKAtjFTh+n0YF5pXJxEV
yZgLr/Bhth/1qDCOiWZfnsAksl5rG/czQCHAGI3xG6eEZRpH/TXdLTvZCl3E3aiV
FJqQDyeW2oKKt/OxKldFiFsbgVj6d4D4OkuP7osajBERhUW+TpX0PJ6oWPzo1UcR
xEOOJR9QaonJBYI5h5gaXPZWICx182c7yQK8rFygRSG+YuZe/TQNiroh8GEEutNa
1yo18YtTxcC26J7SAToLkQT5KbiAozVJrZsH3GxDET2PsJPSQd9tO57JjlCLZKcD
9nXIa9XPazTnRvAz10Wj8OCccIJrRyYlLFzy4x4Dt7TdpM8XcTVR50J71dsf5bDF
F6XRVJlIlw09Xfx+bN25wtnLCx+K5r3uSDooUc4bUl2TDuNbAIDihn4Q4WfgWb3I
mVzUeYAwYNZuwSvsHuROSx+/KJ/IqirnH9fBQXaiuS36CDxSiBOA7gmpub0EVAcg
wzjEWUrVZL0/pvekS3k12XkFe82jwfSK5D1ZCUw1VF+YOLZS+5J5evCWfHjotJ7b
/gtJ5hvYk1GLPVnVuRoNMUV87ZMhGU1JFehAQMhIPaA8N/QfDwj3Agqlpta/jt5D
sfbnWwAhtGvRqnybFQy8JwtSdml+EobCwCxF8rmo+czXrCVEzqC/qd3j4IphOMbk
XWpJli4M2kCW8bN+qhXkTKc7UWpW2iSMrPkzEbjzw3nxcj91qGMzqxGH8Iu5kbYm
W1+Q9kNr2zafjPLA3ltqpfcHGFPRPCYUALIQStIFXPDtuhQ5MxFFc3YKcEoy719R
aOk4X8pSVnK5lCPMSICo7atJo1IEu7YIuqYTq6kttOTEPdZhPtuaX5y3qeJBDu/s
vnsa6WarOxqdmjOWWr1wwik7sDB8a+Vg3xmJ15vZh0A5lAc5+romMlrCxkTq3IzQ
yEhXOIBwJ5yaEtyP42S5P0zogCxyrOueRDgwRSRF3N4l8QxK7lCaUEBTAz0EeqD2
v3zWRcQmniAxk5RjyRdDJaBUG0xPezQyAkm4WJ+C71utZRuqLY4YFbzhws6F3glG
2z8Cw7QbV6pX/O9hRxRNOVfS3PqzvJlr8exQghBiDOdnRs3EmrwPlIpm+pe877E+
Vx1fUwyeUfK3bifj52BpvSLj8A4buUG/dcBA5Z0rTI0PEXDVmEXG6sPeqoy/RV8q
dtDrNGcdgKW075GQt3XgxiT9J/l7aBbY5QfbevLZXHo3RRFQc+XzRvMj3i7Uh/U9
7s7tKNpaTOreEXicZLIVWI8FI7NTwZ9nWbU5H1TJvBZ0phgh8w1uXmwkY5xEsE2V
SSumyOwF2CeDSDTAVTrCIHXqnswlTCkYAB/nCZU4cfJRRXtWjRf1PIie6RPJlYPG
m8/ODKg04vcP3Y4Z1Sup24ETSsl/bU54LNoqa4uLszMy3LbXk/+8VYU8SoPk5K6X
zZznudBZCRZIBc0S3S5PSN3QOACWQsU/dLgGFdYru/7XywmLvyITuDvMAvljlo0s
BAb4k+Fun1IYCCq8npykgJrzGnbKzTZ7FxXemv752tgIv3LJdHCd6AvOhuLVW5A/
bC0tnEdaX/MjErNpjuPxe5O1CbzVwxmbjzoxvf1RyP3zWh2O+jK4L+HpyiiyflWq
hNglH4Y41hWLZZWuG+KKyPa+y4MStuoEmVtwMn7JLLLr90xS48Lnf4YgNDwxtvOY
0YJMs+jUHlc66qgjDwyI+S9B1gbd06z7qGA76BFvtBRePcBu07XugtMw6P4L/7nQ
I6P6Ity5G18jnvAulzoISFOsedev8CBXWVBSSYR/ccjB3QXohqJtuGG1gyrUs/SF
d/wNRj9h4wgiwq2zIcjeiyd5iTnMh9UQI3+JVBYTmAuM3vNnF4kmpzmfoSkizTY8
g4zNIwtgMcV58UNCos5NaiyhxbHn9WDrrCcc1UqrIXDxpHxYc5XfQXqMXQnQzaeR
XQQzzJ9w42r+ohOZbwKxMpxTglvoHIOfdv/6hlMIceO3XU6NMqhqm6QAdzQuO3q4
e80DHec+p3bNzZ6LKlgWfkRxm1vNFnGTyq/aeYNbel4znDfc89NPIrH7qcdSEIpn
6WEZBxFFaW/oVLv4IRfhK5o9FLvcXtvEh7i5vTEy7dw5xMOZA/AJmWQC+HrC/Bok
JLoxGFRUO9N9NtVPBW/Hbi0EkzDnl04sETTo+l3C5Hftl/B0lHdh9+dcT6Ywp6qF
ujalXG8D2ZuPTxs1DTYJWGtHC5fKtkWRMLsaSIylqKiwztuLIPy6+lY05QLCcKrZ
G/Yvizo9jz0h7R2TMbNJHDwJz1psW8b7Yj06pfKkznKZmLrzfFvKtgQ3hwXcSf91
GPjkI4p1KbG2Oq1UEEt9gk0oHvef2vk6se246S7uwr2KkN3eDhPIIiEVTXYHtk9f
SZ7Cl2CRK5cMvmU1Ny4ykZzza9nkK8VZiU30HZPt6OwRCj/d4MCHQB49GNMurS4d
TFRjqek7ongf0qceJvdmNjwXhyQd+Y5SKPhfIUBysFvjEBDLDaQ/RI8kCubtnrbt
ZPtm35ipAjA6ekygMHx3ONao0uK3ArxmJdeOlyKJvF8m9BVWifawRn2TB5c2mgy0
oGOoj7pT/CP8SlzJ8exzWwcnKCn85LgsPARam3gmHxku+Ln/mDlzzkXzfX/IjAW+
DIPluUKNgFe1KyMQb8nw8KpYfybJ6pmkLEhwZiWOjB2VuivUpY3YULspv5eL3dzc
dmYwQt/1mQGfR/LJ1GI6w5ZlxEtwI4GPeDG99/EOuG3lhCF4sWDuAsV9BERrS3Uy
haHJpIIHml7gxHbsTpwHtY0s4rRseW4bbpluArFFg0smpmfAQfARsWXX1s/d0bNS
mfb7NigfTh28zfsx9C/+jDePrwQVwHzVLW3WHZ1LqgCZoZOlyHoI3bPImdCbbA5M
/50YYxE0sEfTEaqNRZAO/GJUPgr5DbVjcUEaM3SPOvPQK3A1LWXL45HXmMxrcb6g
H3TZhbvguC9MNccFVW5pPK7c8RK+NzHDVtEZ6QrmdGy6nsvAtCNvoVTI4uu8tyhk
qNxq/dzwLanMVc7ofHRdhGXInTVdh12+2mULSI4IkS5FoAGNdd4RADRkSG91Vpkr
gaeZaM533o84C/Wz1QYHSUzKvdQf6onyG8qw4kh/AU2zZqkCOF+0E5TrGydJKpFD
vzjojgR6QrBs8Z8pMv/61eq+rLNz1s009OXYxaTvPGh39unkg/rgonTn1c2onuhf
IRlTf7IpmQGAAZuypP0XRyiegSevuJ0IbFqOFdUO8zBWwAACqWGR0zH2CfBTGtWn
1oM5qJ+3BgY4VqOEMAUIfIeHLTy0AHEjOE0Xh8yVUdkN3OccMQI/Ex0KthKihIQc
la89/2TBFrDa2KDA4lpypaiUZ7NFMUWlWOqtoBf2pIakQYGR7uF3h06Gro5waEsU
Qfvcl7O4+jemxCDZX9IRj3bItWRJokJHbDJgWfNbAzhCG7MnRJtE148Qmv5/V6kx
gdVXEJ1jtqsOpe4wP96kpM2dNhykR7+/AE94Q2IPoe5bbPo4iLl24VdSQF4/2TRL
wUH1q3GbCU52VzfqLtp7zeE0axkpZVHXw1sM44tungoxw731/EMtxSl9a3UvMAg3
AMiJiwJdpbd9iWf5l9H5+jgVG6A4kGLgmMRud1UeOOlCrDJLLMRbisco4CSZhvu8
/b0wRqXrEbAFwMUNr46WeokW32T5FouCWiHiNKDrqN2kdpflnIWa1xCP29Kh8xnU
8ZxbIpn9pzo0D8sFZw8k1gWkoHYNyow19c7ekrY3oa03FQJ1GBAv1UkDQ2Qv9UDc
Css5Ea9jRZ+RelbmKNZDxOLRCn9ftLImnG7g7TDfc7dytOQcTPYdTFwW/s6AeZmP
2feseLqIHz7VCGctA+zaDk17z6kLy598OllaDQfAdzjwQnhmqtGImUqbFXkpZz54
qdFHuT5jw/FJbOkx+zQ8HmcRfqSJYNhkXWjCDKXgPFzLVRtf7NpJU6/cvdtReKAF
dXj7s7S6X27NXH68TXmct4YY+X8mjOGO/uy3O34jqfIyhWKaH5jvXLtjR4IopLxT
A2nhTLRwEgMaVsPcfxV3DyI0fIyTDt3crGeYq1vwQ8PIHvQ23U9ETK6ZIHeh/aWU
2QNc3mCh7HLq32Dx78BqI8AC0r4psoZfiacjUtrCja3On43CT7u4xI4KZwg3pB1E
y8aCxw620XZ3pkNxGNzpcEczURW0W8jPdp/8h8nXRt54uRcmoAalKbEzuSCfXQXa
IMMnKcN2sqKy1J4Xs1Tog1qxPabr6rCdqSea18mXm7rIPaz1heis9lmmYXfbWZZk
wda6K+79OsgzIjUxBvYGTcVRtJJ/6d8hrZa294ZxZgoljcwbghBE+SKkiPYBRXj9
91pfm5SWJL543C3RHur727XN8flRzBUg+JTugYfxryIEM6dV/h/mO5qbzN2F+ziW
PgOEZvmgDgHARzCzSum87uQEhKU60KJZ/QVXRRUhOvYAfLsjXbVPbvdoRbOR4SuU
Ai5qK7MVPRWX0gwVz3nIYiH3C8IkeJ2/2PYgUR/3wLVjmdtiR1oElq4VCfC4YoI7
4Imcpcti0wZyVzZHRmDwGF43UQdLi6Y9jPZDtttpwALEhQaDsRoVUiEsEofJEkr1
dBT9sLkoOcWh/oXSbBgIIa8/1z/VWpEXjo0iPu67XKG5m4YwxJkBrpJccvXnpRi3
O5XwMNotz3jRHSe/H4XhC1nRK9Y8JJUbWFANnCgev/0rwgkuZJ3cEZSSRnM0N2xa
VutdwuoNapkg8xDVBJBi7+5jKqq3ZfIC/68boffCcas2lxu0phCQnXPFkQHidWK/
USn//tAGBWsggMyqpjxwgID8umuNpUFg/ISYwnS5vRwDawR216YwbKA/UH+hB3uo
y+ukkoJmD5hsM08OowLL0g2jdeEKtgNo3TKYhgvFSF2neknq/+0N4Rt3KfWI0plz
P+Jm7+qcSgkbwAej0MSNNioAOgcd3qkQA2i/1zZ6g2BTTu9SiDzAOipViehgCFj2
PaUvS6c5GxWiphzJfGDDDWLBJJ7WHyuehHVc495P2tnCpiOIFUEQ8EUj/CrhDAjA
0TMfqV9Ys3UWp+M9WIBegy4E5ghTxT1t8igElMr9CMWHxTdGGMh+QylTjwQHBiQ0
TI8w1mUY8+BaLrqfr7X+65SBsvcbsSfAtAXnMFl3ThEpYFCcygVlSjnjrLeHnkT2
Q/kZYuOlA0oJo+iiiUqrIFP9Qiq0lN53qp+SpAIYRjM64XiNJcyCu7Sef2tP36be
B/FpGgTrU9lG1+0O6jnP4/Wc9BfQ7l7xHMduRjEcpb0X1IVTDRGHEQzLhswotOq6
NoCMokCGO7B4jO39IIoTTXq1YANO9sl/qlde73qUpW4xC+q71dhHDV9PUJgXcSK2
xKnNKp/eZJLkjt0G/JI3Bon988Doywpm5Ki/qKVOUEgPHNz/ucpJHibZubcEyoul
8krxEpS4L1CzJZhn1offoNy6id9+tTu/mCbPxXTFThIlJYP3swejYquJpqh9MtZy
qa9xze3Ln6NP4YmfkddRWgqw5oFfKY3k1pHxdYyhX9R9R/U/w/Yl9K/sd1ftkXky
9m569agLgq6K5W1A6uywFoOtJRexOOjRv7gELGbkBk6KtadachWJDCQ3SNo37Wek
eP0M4XgmwUiG7e5LyMN4l/OcTLu9evQslpLDAHmmsnf/8452BCqOGIpAg1mrvy1V
P0Mmx1uJN6jvyc+LIpSSHZnGk4aIqAmbNObSNaFQQTh+5tJiEn07gGqbDk7K8K0E
c7Cx+psmfiUyuugYfRpSLYw2keRSIum1dh0Jx8Zx6ptIFT88LOtmDnjcq7dbrGt5
u79BP7rq+IYLeA0kmKEDhxD2llos9b84AN6Tmyjwk5zhtK7BX6YtWs50cAp2MGfp
fo3mLB0rvtZ3i24OBa6EYKa5Giug3AFTU0rFefdd/XUe0XWxxdBOrAx+kH2ce0sB
qEp8ELnufgQ3Qo3osh9txefjZO9riJv/PpKgW+P+eAzRGWIJOerwiJ/YUxiPOaiA
hgiKaTrthsRuyHY0HUl2rtbYgqfp2KhW2UX/D46wiEbYjU0OsUuUywCnI+iqS6xd
ppOvbUIs8jc4Rfv7ZB3s5Kr1RH1y+k1YF9/4aigaarjbMlRxyFGgV9ZjB+iKGBdN
l3tzPuh8Z/8KwyAuuWGOV55kKvConZdiNF3QIHG2f6huIiaGjH7sdmMEgxUVDzd6
8MPjGDGvCLccD0XXi6/W1s4w5tsQMijfU9WP1PTVRHVadGT7npE9xrqUZwvY+VF4
pJR/1wU45oZhBuX19rysCBUPRa3RRTb81x9fzIEiWwFR2Lnao14hVU89PxeX4ePC
aErMm/DGsIgRsqHkSpz/TnTkEbfUffOYZUUuqXqK3u/ZRPfUfaTac4J0/P/zHZnt
bI3S5ykPFd3o8dK1fhATdZzbcltRlYpzqZ1dUDmHSZZBAMlf2yYxGKDcZrjTAbx+
Zoiss6gfFu+M5NJr+E+PvvwnRrVYXKD6aoz0o+oxueCM/J+8gV9aeeoyesnSw3xI
hl8+eoLsvxDIt88k8YTurjb3qpFHf+UFq9Sj8lEjGhoxhphdfjUf4WfrHpJzsA8m
TFRFSgWEWzzr8MDixaHNAEv8xaoBVZHSpBDf9aQtQb9aWTD8yRT2uUBknutaDMLi
8VEg4Y1SVOeQZ+KxaDK7souh8Amg2SbK2GcYLer1maYW9I+2JDFfjzv/lOU3fElr
kul2Yk3oocRS+5Vh90gSDrIg6kNT4acQkjcbsv+OI77Mpr0xFcpUxPF4wIzfHYfR
szb8VBumRCMUBVvRWexpPtIMvrvf+e4lx61VNOMWJIX5hCTKS82O633Kcc1Q0GU2
JpLQ0E2tUY452dS1u345+tSMjHW7BHdFI8YKPT9IH6sFzZv5vSsSMQFyKzyiOiXB
jJlNwWwEZuIvMq7fEJeHqkAHKRjYYHgF4giVEi42roaJ/VomxtUOXB6ZR/WWRJcI
HGVa0PocSno9izroLHiH09cUz2+Nkg1ztGCNOZPJC82QtuYbKlu8xeVG4abG+y/H
EL3sc7lchFeNZSKp7VC6zoqPk4Mc6d/WEg/O5MDjK9Gg5tGDxl8tAyeVzjd3nntx
mdqEVCNLw0CT9dWySNgYQkn0jnChwh+ZxGVwqehmdIbajYuoKSXj3++RZam+Fv4I
CfPgarsfHKZvjzhqpIZZvbz64nBP8rsMf1VmJ/IRRIZSK/uC8Ul+jGpHn68bvWpb
VcRzIbfY1Vu2HVa6MByBtrOa7JpuQaFhNhCto2okQQ9w5opKe0iV3a0CmnbGgwCF
mr43FsKXxV66L8wiDsT8uCiYNhNu7Lvma8lwetfan+Mgc2PBSeD9VeHMlH3kGXL2
d5FWqqItsqSqy0nSFvQxYy0ny/EwUf7NclCMeW9F+LNQrLS/lCifOzXzSVWftzIU
DteXm3scUuD5eRHw3UAoVOY+jXT8zKNUQ+a/nEfxwZEchlRoybgJX5lltetLpZAo
4zy3hX584DIMATTxlq9MRck5RWpsNBINbwT9LTEsbAF/8M6LnCvNc6mYTdpd4TfP
y+6OO9/GH+ev3fB0fgcDZcxmMnrgRgHV8VcSQ3xHsCjplFpyO51jH9YO/Hjev01C
eDwkDi4NZ0ysEY7M5UYzDows60uOmI8w8AbU2spB7esP9kqYGBIwStUhwVL18hkA
pif3qysLKNRAtnqyJ3Tj7gNGRChLCR+2qeNKgtFs2N2bNWKi9zjyx8b1Vd5zxBD8
MzGKvhT0b0OaVd3UapQjA3lGAOzj5XVQclm/hY6xI33pZaa1H8XhETtExujEuhdB
yokR3n6skVV79yzDdmfoUMBRUMoid8CWY1ldQeywBlL7PcM8K7Wn4CUPA1191HK4
zNO0ErmVs8C6sVbm0ciMPVwXqSwrEnuSL3Y8OVJ28UWSCVCMVRlufukFmCeZmWzT
oIMQQLG808/HWSoq0lgzuaEyNgz8/Colh0jYM0Lic87456VXHL6tnps5egS7dBBA
k9ZHrIhORF62eLHPsMIKh+ACFbzElJB6uJIvdY2RHmly3wr+XdnmQAc42cDTfGJA
p3lznf8+HfhMv9yfxVyllc0NAE2tdlNhyZuwgiX6hO3Acn6O6RK6kIErTUijOvk+
7fioV4le7m701xHJJ7dIzeMicVYUfsxC3n4b3AirI0jJXC6eMiSzBQLVrs6JKx9+
klH/aNp+pLUBxPB8c3fNZlu7NHX+CnjtCfmm9RSc15u1/s8aEnmau36/tUsH9mFg
ZS7CIjLL69LTXKMB5f7fSJYTElPgTdjXwLATgTPy8oLu2ls8ClzYTI5aU/Wbrrue
6rBVm/mZ4ah5a3Yf8Swr3w++zOa+TuWlNFC8In9VsE0JCCi5EdbKfLVtAcsvbyf4
TTuC4QGaFaf1aSI/Ef4Gyfq1HgORRr0UPBc0tCrlE6V9zN7it7nSDWJn6/mWtXy9
wX8GG0i4oVc3VcG+F8jt6m4nSZAmwWJuvjiXyHA/Yd2FWok25cGjRxHrxsMxp83c
l1xCVd6juOhISgnUiKmutKuLH5n7gFWAfh/hOuHLJcyFAVvqkWk7S+zhlmwevC40
z5ce7iU1fA8GxJElqcHSZvZPXl5ncsqTUO0VTlyp4I9dcWtQADVsJFZKu1OjkN5R
c3bc8AfKX7tby2/TJVGVNKD2T+ofDEi1K41p17Gru9jvz3bwgRvSbalbuNLoJ425
hW11q3Wnd5ptxgSL3rpsVQ1rtTruKY3qux9fiWVtXaY573L7MNkpkSoZ34gjvaKB
YUHc5o0Sxn0RcJMXwQlqdTJlKHGnwYQ3yiGySRAEUTeOTOYZSu65r/IRmOmtU74P
TlJ+5/vfewUEfX0pwfRbK1bQO/jcl0p+JcLYVuw97SOhjsvf8Im+aJgxvacm11fJ
dVltRTKpzFbSAYIrG7aUHDCkAVTEXRfcXklq80r5nAEZHtEfuDZ/5rzIFcAhU4tB
OqUjkXGIJ9abEacRcFGgyduLnx5Kr2rV2Vzzgwjn6uPgkneOW1GdevKoJYwrkaRL
+xMi8g2i0E6Jt2fd6rFbPiYXGwp6hqGFHIyKKS6pr0QiUZkMr9tZmeuLjrl3F8Mg
gfMbEbB0ghEQ6F77KS3ZN0TwVW5IAwsVFwvxxGxNhNrOzQyGt7gZvBAPBPxy8mJA
IiwWoX3OYQsdvuHeTe+UBrvZfBR/ve+6as5mVKCO23uzCF/ys7nwIc4XYTk0KdT/
oapAlkscDcTg3jbOykHCzJuYxKMN1IVcjp39bsxkicwOwGJUWzI7RuLjSsSEK6lU
M3Cn67Q9jdbOa+48i6F9YlosoVp/OuaMn0RluZ4LT8tffkssppXPKUo9W9TS9ThR
npxiG5RwlN4v2qe/u6K+nhfgVpkKvhXGlkA65BqEX/OlHcPBsdT8iXuTF7plVqXJ
T6yY8o9QGNA3wPRiAowefGzL30cTlZr3VGiwHQVRNCSnQrv3RCcp+MJQR7p4zT26
Eqo2zmld5X/c3BPRIPP8YkPC+9W3BhaqHMpyHiGbA4hYP5Uq76rYgxgHWqOFTs5P
JiqPI9ZJkgkBqKpawZ5IQCsM+1/RdhpGzxkaeKydrGx4pQe/rfdwqZOfqVH/Tk9I
OKvV+UWFKEOp4/TMRRkuwl04wv4w2XkW3pDVLdQxu4H3k6h9aG6UCpoYF+4+enSQ
PJjGzAdTJE3IZ6+w5z9IMoPHkIvbQyHM6bYCnF2WR+pu+M+YdUkaLE4Z37u8AG2e
uUlVwXQBu+rzUMAwt++8IpmHXy7HtlVynNAwKUag84ZwX/8TNMspmW4jR+h0jYdK
7NXXPDUph38qgOr4IC40/SYr6Yme1b4J7ZESQtsy8Sjxt7DW+nmIgVEYXSh5wpUD
siRftxbsaQ1dJMefVd645RSL5a2Pt3gX4TWTpxG6+A1Z9RoIbNSv/Rjylg/iDW3V
HUokTdiXCg39VcDdxvHGos37rszflc7YviMUsRDxLsB/BQOHtnTce2AsOw40bhN3
grBwPe1QoEVllcgswNX1wBIBh2JXcwtJj/11PSioy9mpczIxhnMKFJvGpnthct7y
3CBjGIhy0K95PqU30iWQIVHO9nGwjBXh/z6+P57ydTEypshM7PmalkotRkf8Nw0R
JwPjQnr1UChUdgjZr0aNaiGYW0JU7rtqCoYRdQVMkPBWnaHm+rD3J/Qp3SxspUDc
OCvRAAoQLnHfdcZWKrsAOa/oY79l4aJlXTJ+//FKxKKKfCfqhl0USgPVmi0R7las
coAsK03auncLaT9GrNJCEYh+jQejh1kHvzagqbJAa+tAi1Sloe3kkKet5Y1SCxzN
zRF/fw94t7CCeMQ+fxcdlz7EfDJWspFlVeAMnegCYfk3CWTiAnAjHUxYxAdcGVky
FWDHG4zZbUkC24UaDG/6YuXRBRWkYMQzpAhNFIKuShp0IT39MZ5zv+UIOw1jY4MM
8RWurcEutrp01vopw5Q4UsZsGvRdPtnjn4DZ1oCsELkAjuBqJ2rOMgYlTEeAoYHO
oRkvdFzMtU1C7/PA7eNXooNixD3lqsfVUd8aNsWtKATUdabOMDfamusNdBwvGt/C
OLIcoToWfBma+LZpZBIAp3TgkPAwNAl4CLzLArnbKNd9nGG5ZLyzBc+qpxGm4mwl
DFxN/bCYnG8a0mNYaEVO4KlBF+gpceDhibXbaI151LXxTq22EDsVtLVOczjGCy/H
lYfaibXj4b0LmqVfwUkNdIgU1QRXDi7EA9kU+VD6OCoUdiN0EEXGPuni6aNgR9sU
KZWeNzNRKOz7E9xKWvjuvvKfNWLfUti/r/p1A6pnDqI6ScjvdgGxzo9aaOZ9p98v
u1o6FcYQvEANZ3ymIv031L6ohAhHL5OpzfvWOE6vLze3cjcDBYptXXFmpa63QStq
k7AKF57lnR+GgUQgYLA9kD8oU+dctWg+78hQ4Sc1jomztjXYRFwClNR1VA9cEEAX
t4UKJlnyt5tFL2i+b0fgHDGybSUsbvCrrn1U+iEuBi7/39v0ORJUNz64xOVEN/99
F4CxBVCodNX4RpwUg5g4HzGsEy8KHKDGSKUr14rXOj2AAOcopWE+AKs0lI1IaWHx
3Lbn9qCEi2q4UICD7+LZAkp2on2LdzBJYt8TBG5rIBVfhzxdIGqCr3pnihBCuifQ
6GV13ITpZ7DV1aNfiHc7iG8u0ORaWlI+d9QC/19fN9/co2mJ3SbPYJiuKDmK8R8A
dNg0Hi9FxPkyhqVuDZcjUsDk/0e9IJzON2Lihq8AEcPwJnsy0VSUv+7APYoklAjH
nlVOPS4leKEPGSpS/UILXfWrPajADaR2R4/qJr/e4Bz23TPqu2pbvh5L4jXQxvQg
gpJhbE7HlOOnpO6yp55PNNRdsvt95Ylb4fvmTkSHrEIFXrlaQTGqkjQ7vedLSN7N
0ZiHe2jskFYBEwV8gxQMP6VZdzCES7cF2Cm6DHqsiDVbHArq+HTPGx7bJ2s4kWcQ
+rHQhKgMCXd5GBfZCNUEpyVrr2JE6LPwrYNCpI6NsVuPtARI+mrBDk46kehYKxCw
XuQUgOTZiymfNPbJa4NzLr4A8PaNYw6B3csIfoXOiIs1k7kq+q2/x7Xo4rsLJs5j
C7MNN1zX6o6f93KDZxp2VQGSwg9sIxG9zRJAUeOz2eg0+Zh7fQHeZqO6xxJ3ETOF
FW+pKy/uFMaAK6yBJJuskCXjhQZs6G/oTeDloEbm6RbTAT1ML5dSAOaXIjurVUAv
uX+CdBLC0GZNvGbqJ5m/iSL4K41DWEf5JPxvFkZKcBA2bGAOxRObCoiVmnOGuEMQ
qbLS+qsMtbR0Pd6+ToCh2TQDUeiw/543Ed5vBO7h2OtHv1XOF1Z4RSvrOZ/w6sL/
tzQ6bjLXxhM04ufU2I5EBXukS60n9C2EHluaOMHAG6sOtaDDundPVUrNHxuf8pZm
rkBwA3flw0d+Kt4I/9SeKYUKdduqf0FxTNTdSRv92ZcXDa9hO/nSEc1/+zr0RZbp
HYd8n9F3N/QJXvZNcGMMdNHqVAj66OjXCS6Oa8cqdKNpUyAFrzMWfAZu5Z5Ld/rk
cXxx+U9I9ud+fEIAXKie3CisTHvrJR6dfmHxq/EIczmZZ8wfQYmzcaycouF2fMtm
Fs2cH59mw9giYaPjMk7NhAxisd59wHPiEqs0mte0JEj7mnx0cJe7MxMXtbFnM8Du
03Gio1ooUiG0qF1SRKk5Kstel29XpIuYvVGV0owscXzJA3h2zox1qRZwQdFsfbjP
r9a5zzrXjVK/4jwVTlFF30CQ71OyWZgLUzPxZiK92OHU7ldSk5fQ9dR9nDJ4/jOR
QEyjw1jCXzCR/5Mg/ZGMENYl2uAi+u+36oQad4T6cuMu+frocfGtys4+qOQlL7XL
sJPnqwlkvlJfg5FjJFNJeegZDNRsQpvovHmSm4w5MqIfxri7yHLdiWg6xRtWl1ly
pxPJDrAvaaB2kGbdfjSDQrFhWNup5Oh9v1H6aSS17q3Td7u7Hgc0Tv4q5LN1W161
2OS+2R7N9oz6KZkCGLNCB2wYGIFiFMPzNExwfFYGe3jhdvTIZ/JGD/RP2xS/Vn7K
vrL+lYvD+6YaAuWZpUEuzLx99zTuGiWJ2NCFebmJ1cSTSBa0AVeotEuOIG46Mbgg
NUeA5GSxGsdvGXLDmCdTC1XXcE23yUbbjTbS4bjP5nJvf/0Q4705fr9KQn/zbuZv
MjEz5LXUq/0yKJkTrWR7nhU3nftPXA3fYmosyonNp4BmTIYSY3NsFJS9n8oSKIVD
ReWd8ZirJJpkVhFNjTVwCknlabC/VA5Z+3Mqge+Q/H21WhwJYNR4oZmmFTcfuNuF
Wwbj5SrohUK6t1oIIqw+KcRytZrrcFKwFvfN73t4QJtHnEZKiKzhgpWqJAm8q5J9
gqcI39PdKqKxOY2ZSBbsmyi4sN47uB4ACyoCsbd/iMTb9aRCQHo/W8yVyx+DCHzm
spkAWJzBKl+hEe020ddl5NmQzffiPbMv4u5mkc6leNMb1n3gAtkhIH+34doJuOU1
Z8gS7zbf1YULZBcyYExZ06z+PDQfyfqwmUmplm30SIEBF22WO5qkZWjM+yzJEHqM
xyNh1tgto43uwSYd2cGM/5WHuqmVfxzxVL5B6DKpBrL2UaFNmYlU9j4dUYhC2VLU
6q0OZHGNuexYpUFkN1j4isMMFhsVK023TeJ1OHle4OSVIT+f8g0AxYdorgLuR405
W1tlMdDg92+10tyX4bA+qEKAip+N5q5YCmDumDDHhiEBKkPV9x6FjaUke+jcTMDH
XVw5howF80fz1Zy+jOySLkeoYTROKHJAsua7hAH4OOdlOEywKS5dHRVPHlJlSWyB
KFh2hM8+isFK6Vkd8cQ48X//7CF8Wu8PBjOZfs3Bv4Q4MbDFIFPppIUE7c+uHQiS
BdcIubVThlsGVzC1d/YSp4Q32eTW3LWhwoKdPq92ODLx0JIeCiWZSpBIPP0vDE+o
bFufpPpxLHQyTrbmhP6m7w/VwdRFYWJwO29r0tYqrM16dGuct9FxCPnCPnl+4ZFy
Nza0aaNMS9whszaCcV8WkuQr9nYOWZAmk60AjiQ1meRp9QwzhN9rGAZtylvFUYHh
/T4GU4zDEw410gvqGS63PQ7mtXp/ClB35wvXTxDahaXFFMnzrfZXT9zlLgm/tyia
uJ0YyO1TDPs9+PkW8rLUpVdB2BgJNixPyL9RpURfc26mwcLUrpSIH8CnpYU+owiy
0MvXp8j4V/sSEAgMoyC+t2BQWqH23+kBanS5WYFPl5OKKU/Xt/GoW+8/sPIXQfBZ
AxE3ec5mUPejDG3vUzDqcbx5RRU0effvGG5wy9bBZg/MhzYAvNZpONNW0ZO+LZMA
tydl4ZMxLMptvSzxS/ekFIAjMk+SshSiRYlW0nNam+h/arI0cHhi0C2sySrtCRxU
/KKP+Giqcgf+x0at9+k0BsCeR91nTzTkR3yo/kZutT+uOGb9H9EE7slXRwxWQ60C
R9QX+BnaPucO1Ag2FuNrizm5fY5aSGmm886dyMtlmTA9chjec2k1ASF8hvRQ8jJO
wYWjGw+iVO1++g+SoQiSTcIdfvvwKt6OKrf1IdGpG9ki1WzRB8DCUsx1XwxiWN+1
mBkmyW0rJBlhzXU2lyaRKBxZ3L26VCWP3TfS2F4l1ie3l5kvI9GOfQXelt5SDzuB
rToAgsotMrnj7ELHeSQYv3/aCUNSq28l9OLnkiKkZr3IsDKJ4eJxiJvqCzHLkI3P
tcInQMR27a/bRC23OSLRJlDKukG6HqVqr6gsGmr/aPWwZBZxOLvmnEpaGSvorE2L
ShPDSDNUPDGe63755w4czd/j8EyQP0jiYaMsjy98b0OtxKy81KiV64spXBwNHQyY
RWvyud3tey5hwBlD2fHWMZyxYt2eG5H3EmvJKGFVYRp7oDoyLvRCUo2fk0bZePoG
ujGrqn1V9rnEk5Uj/zbDPKpTtnSLk/ZPAzsyHg1e01JhaQRgZQkYl1sRM059ZPvj
GLd5w1LB1vPAINS4dg2aD8bPfFVytuUGxhuY64/p3oPnfOpA67KkmE7kYJiies87
t0sQf1Kep9Ofz/1QkpTgw1Y0m/HNj2/Y1lOMPF5cAN3GI2rVZ+Apjfag754X54eB
0zU2to4CRhqWN4rXpGTMIwU+l+ASJeOINas8WbjJNFWgPXyi8bqQ7MS/I4SxDxzZ
LejOpLm5o9oFVe13fPWoSKOultMguIdYwgzZB7On6WeEnhRCEM1Nx5VyrLOHu3jv
Eqgo6GNxNQO4Y1/b58JnGLnjnZ7qAiXnqkru4gwZCi1gVSDOMl/fsXNjz5qdupk3
+tQWhtNF6j1wqnLKMdq7qr3Qx+HUzcHj6DSp8l3mHbPV6oTbRL92pIA9Rj9COs94
5L67oHhgGCVB0oBN0Aq/iBnih3F+YHxo/ejmJy7Yhv5Y7jOIo6pF/xXNGEAAJNvg
dNGo7bL2RwxeEBMIwqNFPmGbG7BE56Sl9ndRjUm5/6FbBdCJR28nhAJ5eJNmjfwm
LA1RV8xEtSIEhQg2kx34OYFukI0Eb1cvGLy4+pB6oWnd++1Ci0Osw/OmnOFIPkXD
cyB2RWxWgaRvxz/J8gW0K28aZ4cTW13n0ALWlnmrhoOd2xFJwMNutYBbRchklCD7
jIE1Szkt1cA0IWpgBFLVEp4k1ZRBjmkmEXZ7/WC5/N+duLQmUxplMe+6OcIFbNvV
Nsg/OjULqLgo1tFIOBGeh9T1WhOR5O5eBHBv+JrUnXCO97zMIweKWHO8yxqQWdKr
LEEtlKEzBi2WneOL+kYTHuInyL0yYmKx0DxiwxxW/wyj8BL2QQf/XO0XDModuoXc
H8UHnMpvOHdxQ7J1ahTeBZHXzkC9m2AZhc3SKA7T9sn3/gHt7RceA57TSE4piq9r
FZVt5T3JbV7Ayhx7Br/IUWJmIv5JtJlFpR6xdrpidqQIiX3IIIvrWeqTTmtkYyvf
7RnCeUJ4+UyaFXvWr4nRYpAwNe6n2mm6HfaCcoIct1K1rLnStgJcwLh2KHsiUQMc
Jr2hPgkunhm6NPC5EaEhZL3Hr4f86AUYDfv8KQ5jro+IFYnj3szjzQjXnEfdDrPn
j0i6y2Msb+hVa+Px4C1jVKTTN3Q++PuUvs+RBwTWCRGhttrIUo0UGkodpUzApe5v
flpEZ8787vOiae6Qn43B8pCgIozLvK7qA4o/7xzaEgF6TvPfclssy9M0KH+51MIS
z6VNdbZKwzGSoaUwUdT7SHUmCUWDaO0DLXW6fLgIH2J/gsg9lzvm4m7EtAh8Uxvo
MBFUBDCk+tADsRqXhjsdijI2nc7ElrGofyGQlvwq4mclhzgqZOoqIa9WLQwwx9xW
NOZNZnafBOtxBWzDz5N+/R3sysAXgNtMVPTkzlDo7DvGgQ0hD6X42m7zNjyHmJ2q
YKqU9U/gND3Q9L5haLQ024M6zMTmKT9mYSga1Y++p/2MEJc1syR5cXcf0FfLKKrZ
ifbBWvE8TfnuR3rj9pIyMsuySWdXPHXRLZh9PCBTYMTFfyr1b9Eg88ENmj31OKSu
EG9RinpwGX6h1WZz0L0dDBF9v8b8DHDPezaGwgHDBrqAIdwMu5pN2SAnXDUVhEms
KKWgR4SxJdRTx7sAU2B1WmQRqbkJDMMA/ExBKHgZ6H4PEbI4r/CgxOxfiKtSdt6M
CZ4jiHfnG+2ENCcbCRILg8/HJOhRu5VAR/1Eahdyu4pZpk2pQ2lIe4lBdNbQrFhn
R23Gdm2tefGqW8exn7Foa8dDpHH7K4Zhm2J14j2jIZdsnI4ZyawuxWdw409QsJ2W
3JWnrqkNYIa5/uNC4p9M8adYD7karTo2iFzNYb3igcf1RMWaVSD96h50DIXMyLY7
1JV/FOavjsasPsRybb5WquV2Iz7pW/whwhUCxfoFfxPMpq2ui3cwEvepL4C8TAOE
eee0lK/dZR1BLpcmOiWL6P787lH5vmad6x1ECph7/Hb12F96WjS/cXwO/w714QbE
yRGdEa5wZmMelMl0MStXfq0GRK16CMemLAg5dfzk4ciZ3hfD9iC8ldt925NoBBBz
YeGsjF+Li9IPnVNulqiEhNxTgXKedsBtsjeiMOxFhI9iWb9Er8WTRH4ZCSvIgfNi
G+GvHgAYYW5hfFz2lASAJQAAxyU10HfZKV4gC6Gn+9RDsTqdPjq+5plY3r5Wht/+
3RzWnIrzAysO3n57leLyjgIBwjnpyCOaUmGM0/a/fBuNg8G6x8qATwlHyPnR6lVF
8yq89PIhoFoJR3Q2NRMR7AJCo2cTjsroh5cC8W74eOEPVwbAZUFlOvmgr/2rgdad
9Kr6dSgvUFlC1Ff5swA17ix9uuHFSyfMztPv1ULm+4kL1TdMssjTlS5webeQT0E8
EjWbX6v1IHQ64VIeENFuedH4PcbrpeC9ETdyDb/Z7KccCIj+a8IhJU88picDmz7F
1F/bGMO1Zfc/tzIeDGwSB9yYtosAOwe5lN6wxaKlMczUDDQE33rXLMnYuvyw++Bj
7iEz2X/cQCVgQ5bd0FWM+CF3AZfFYWkaUpOwULp9bgAtzreRJvJBT9uXQGmA7RKY
rr432oHkw5FF/ve3TApAU8Ym5G4THBbfq/79mkKEgkSJS+MOC1tTcKZa6ohqKyvi
N2qmEkqbQ4mfom2uZSXxaOrAyH3tOQyD+mTIISXvncz58xjNleHThsRKdn97jVxs
O6dcHJx7Z4BTbTFx6uN9mRBDd1qOMiB53+B5wPVIDyZwMl/Kyx/uM9yHvEfbdCO2
BhCoxmu7zuRJjnq95FKomRozcIvB/+8X8PUDkcFfN2LLSC4ozo9MXKetOFHcz84I
TywlHlldsvV5x2vqcyPjpOUL6hDk7FtYm4HWoanw+sUMk7jHMWhCi+RINyCrZu3e
W2sVpOm2F+Lv0oRoM/Uy3oESaDDpuPE/PEj3mTNoMwM22Jx1u3Dk0Rao2HduWoaJ
yEXGNPha16dVW1TBICtoVA6WrkbB6h/gUM8oMd+I3LOPo7YwNSv5HGgg7wPiFegu
vyJbK10wTEz+Ujzi6YAczD27xymdOcE3q021JdGNC8N0X7B5/EYbSX572xKFF/w0
nSgoCe7gRQrFDQA9CBQv+Ee7nX8fxeEDRVrcigrQIWtBDPdBNrGz7ESbFh+/pF/M
thy2QsNjvDAF8c1RS7BqC/f+oGIBTS41H55p5o7CP9EHhimjFdu6zdjdJOnV5Y0W
fmjWSrp7YXUhBtObUmoLSF/MDR3Tt07JQsh/MTqP7ehJRv9E4SHeUYlImCPXEwFk
8wPKiN/Po4NbDOHJf+2PPuRMFNPPhBb0vPaSGKLlmXQlGy+cV/bjBPemR0yKIrte
UlLNUTHbvRF1iwnKB7AEuHxNTCcdDzDlbPOzY7Aum6ddE3qDedB/4veJI+uFc88u
J73sVL4Aoxr4lEo5wnO2T9vWaUw0Mmp5jK2Van6cfXq8hH0Utgb/52JT811dyRTa
4pj/lHFDEsbvGbJBOPsl4y088oH+73Q/tL0gNZceL0JjxYVU7SNlbOzFut+vQiTX
+rEHIGu/E62kc7KhUHrLEtTtRTRWzTHoycyDxgNRENE9nctzLfr0H/aHGMmi94dl
nHHbT2aROSOjT1A3GMoZnb5q6sBjPZRUl6XU0TdPdZMytjvV99fBxPNgBEXGMeY/
rSJvk4Ra+S2SDIrnUQ8k6ylLSTV4tEfDRoFX0WDfs23y9suMb5txydpBb2SL1MGW
8MncZNu/HU35wcIfTsRi+yq0e3ak1QqUB2++o188h1wcx9xcodZBLUvJSm4Wil4j
v8e8hZ0LUFBXCniDCbNbfFHg9CxTYd/FHbqjEavgrMmJ+vXJsQNaI8S7sK54K+/v
xGghOhgjPr343ASkdo5+Pa90I3Lsw7rUHcRfyH/2xsyYIc7Ff6U3pwSQdNptWx5j
e2l1dazbI/gfLslbQFPAuF17j1I2my5qSHZj0G6T629LWzm7ThLcK23TX5jPKnHM
n/+dIdylpSHy869yubtVfvQmOEuqpBpV8uwOhQ6eFhiZK5kMO/55ynv4pfV3q8kw
7wf96wH80TvqFWdzEygi0w0lK2I4YZUddCpl4BITCFhQaSaPniuNWVatTkp+mh68
9fra3btIXsBY4SmOxUvQItVQhqXUlsXSzCAzv3NvTY5nZZc5OCTsGcGVHhsemUag
LW+CMoY6CJqiNXKFSRLWCE6PhlpBLqFDWq7Rpy2CMKJwputdb3uLkXeESdbpqrm/
L/iySTZqoWjpDsvPp1OG72HPXEETIHpaRsPf9VI/kbYHMKX9xapvHGra9NnFyiFW
RRI5CEixh4v/eeMG10fkFfYy/oDV9gk7mwqXAkMYyuf8mcTFVlzeKGd/SMD9tAAH
aKpKTeja6xRV/hPlnTU/8zhyVw3CnYaTYQhtYcUAV+N2jIC+vjqTU4FeBQuwz0cs
V2odp+qk69IdayrqKxnGGmPc0PlIImbotW9OidGR+FzTY36x48QbfS3UVOGeuTfh
xOi88egZptp6ohAymQpn90AMn2oF/F30XlZ6wGik2YNIA2RxELp05FemKQphTgBI
r44i1cc0ZkLdL/UaMfFklDlny3p+xpK+0mycz3eQzqpyUiorCUNPuu+ywzzrVxI1
5MUAthGZgWYIdYbigSVXIu0PzX0iPKonHrErP+Uyh+/abHcW5AGZdZygsHixvNaJ
DtWmTvDX+/MCwjaAM0FWrVrZhgM3Skj76xHQESbM/RXKGK6ZOB65FSfFmIu6jm9C
L7D+qUY4nPc8oGqxuDyOQ/GnpoRoXLnHkhWPfi6gft4PYuS89PLc1+Wql72IiSoP
lUj11rEmLSJuNlaZ09yUkqCttfKjBla+vjkMd6ClH9LFRRtqFDMG+xNExtnW1iKu
kme3KMkK80JeR0MCT0Q96aodgCTYLCAhAUF4VE+yIuMB871wtlpFFgMOMZY+iMJP
EjDZJ3KEHqWf3qbUnwlJuCJzDkQ/n8KUlobJhUyDFgRoiV9ehSv243Fjpfgu+uWI
8FjbohiXO9UG9rrY9GZZqCoOkBiaP08TtZ3WFMZIQ04B3IAiXGREy84sMAiE6qAw
tXnAxX1T4iaDsrX9aEy/cFHj/J61nl3Ukt0hdy5pP430BZo8+1TipBwNAStPrtik
5uqM60+avTIxWwv8kLMc+R+kxTqF4W59Yjyzmx/xQ7nNwv/MEJsAQbIHN+jahgdr
mclHXdsOThJWgCoo0DvtUPawcfsk7mwlSDo6b+6gwtG9PzvyaVOBwoNICYWYuya7
J+rLYr+pxs0bK+kNlcIAEGRuczcVQd9oq5cNz253RE5qC76Sx2ErfsYC7OVqskG8
xv4F3R+GWg8PB9WZArdi1uGI6XVLHCigXQdrmwmI1j3wCW5TX8pNe7Qy5ILmEvpo
iQphimic5vqfTU8BhfLNBtXjbRHl8gcmKDT19uYxQi+dom5q4T3vdqCwoITDJcNa
Gb9qKjuT6XHA0nC4JUfux1i2qJEg3Z3SChwhii2RVRbzJuWcAeHmx3jUQB0p60oc
JaRx3JNUpa0BnXJ+qDOaUS/PIVedKOeEttZZF0A+W5j1vVr6poekT6n73p7ni74G
YMzCY4wQYNm5gHz5q2CnGWKWjg8KkWn8vdKkMTJJ3FCuRZENYK7tHhQBCOLIcAeZ
UOmvM08KJlFXqqpaUbZJmNz6ffevdz5AF8s5sftE5g68QCqSCSncwOSV2JxAFQxa
ueCDHKcTitj12tKAQsih3Sb3hfBmyIKGm0xpIeYuD2JkorjmnjL28JySfKOTar6e
GdMNKlsjUBiFaRIJf/7R9cQL0T/kKsKVNIp/DNE3r0700hw0YbaaZ+HnOq0KQFf4
4AmEWeFIryFpcXrwLdVnYLDMv9vhglRz36SV/Ld9Xq2xNNfIoKGz9+Sm8GiD61Y6
7S34DNFJcsqGCicA4aLXJT/m+I8/luy6BRvCZ8koEa1ami7PR+VNswudpTRm0jR/
4uL8nGsVgtgUcQuHsKWZQGm1SHgUHsIVALKV+BKngO2YQLl7XtLpFuMfpQ7LocDu
ycGWIf7wIbsCnzHYWOOG5Vj5hz6fhQefjH5FCVDTrF9o3DZJB8OjUxL2kD0z3Q2v
go5+qp8uyq7GtJ7+hqPxGQ==
`pragma protect end_protected
