// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p0sPZ87r3Mq8RyphOJ/WR8mhUPy3MYBC+WoI0+/KvNLpFTwvogQVOZbB2DqhHow/
Qs8VoEo6le1EpHt82M4KKQnDxh/KUdagbDQoPu9/bUf5i90gCQyn+LraQix6N++p
BEO3HUVmvd142zFVwskGXvpnu01yj7r7syipgjD2rQA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 174272)
yyqxaiYN23HMBF20wHMftsCzwh/Tw1PIl6rGDK9/5EiZjt5ojImZWTuUUfAclMu0
UQlOdp2CJc/s6HqeRxBytOANmrtHfAUHd8ltFBz2cdDSPXTlmRkB5WbvTNl5wPk5
Ro1F81JryU5ViyGwX77YkgeLwbMRHHDdf+QGl+szM0PlcFefc1hKB/uHyr+EOZP/
MIR4gyK04A5X2RhXKduUY9xsypI9qe8bC1g2nsFtGWPulKL6gyIxTUITU7xiFC0C
S1J7qjjoM+4miLhx9krGwX0BtuwB25SjEeGQFU/VZtkFbyqt7Qk9KHbfk4LxN8wM
eJLrYec761HFHRLO9D4IDSPWUgRzO16Q9dxo2YWzTXRry+S/wSwOp1J+Ume8s0HG
QpC0lVElbETMgDMEdpLgEX3j53WhMnT8dEYSzPe0E7yReQ4l2123k5eJqRTrfGjG
vAvLQvoNN4/M3jeOJ2kpwchUyUBGSMMpxZRrsqHCXfYAJjC52ea0iNZ7a73PaY+R
nn19wlBkJyPpUTbfH2eXbVoyXrEDHkQ4Mn5FxblB0YII8kgC90rajQ2c+1+SbbBl
1fsR7NXclw792uQMoZnZf0McbIf2GvCm/mPYyP3HbptVIixtOTm82r8L76/jYeV4
ZfYqvo470l4B9ty5owsH1obpiZOZxok80eFuaoT7apNuOZJMCxs6qPt8gCGB9pdf
4jfdmyf8Dk6cjIf5kVWYY/igUuZnbvjPU9h7H2jE3uTtq1sWQbJQBoiBL1tQJOKZ
oGRI8M+fiZ26Tl0vXhc3wvpwEMzgCaI7sK4dW15SN1vY32ZgjmtykDSXQPl0tGcK
mWg7r08laK2VoC+n6LC5hMgLl1xLAE1b8JlBPT5bPPtt5IpjqZgsT9RhMgKC2oSf
eXA/kcWLBYhWaEZ4TPzf9waKZx+I7lG+K2OjCaZELsV0uIDlEkyoJ9OEzGPeQC6Y
86sZ63KtISu+x7jyG3fTjD880p5sV25Zh5pQZPnNH0aGfJn3ZiCqzDnvC2mfEFHR
IpXFz1wY+93fUyYC/6LbFMjWMJlt1ry6Y762vPIzxxQ7xXpqeMPsR+o97LpWL2uJ
SxdW2npxivEXLp2vcYMJZ8Rt9KO93PFAyCfMQL54igvvBfMzCylBIoEIAwyjGDlp
LUsePKh2S7sOZE5TXtqY/Km7hG4oooS5YPxRmauIcrY+hR1YOIBQqg7JCen7XAOy
9H9RAvPajfD9xiMnWjqDr5ZpC/e1wgvzVu0xgouw2GgKzoXibW/bDSM4Rm2X/hJl
OLnWr2yXwBEBhQt/2glnfUJYRdXl98XFx1rymo8iGv6YeTZJrtOOaVoJTIOXIlZQ
IfQRv/y+4QFQH3VlHjUyx+kovp6BV2+ixLn1NQ42lbtnjZ+DM3sauUDiBup71jAO
/Q8nZ+9vXziUc3rOxqMXR6QbXzFSVLYEzujiB/GWQ2I+e0XDhm0+3rsvC5r/03nN
q0e8MjhKngcEZaavgyRrwCzu6/zkDXyVJZp2gn+gpv87eVexFJzC/h3aIG695LUm
LRvw+FF/uhTef+dv+fIEBI1Dg1Dc8NGhy/vdNwXoQRMRZaKXDnjAE5GVbFDCiCt4
FBnqDgepW+64aJs+JvgeMNP68lBLBGKu9iSOtaN06NWOI9c8vZpFwrewHO1Ayt10
P4t1bIT85SuQio9LnZFQT+lF7gKgl11VDVjp4da0bY/2vs0gtf/3omkVE0EYPUst
wYYpXtK/sFmmjwCZtqNUZbn64/M0M9uVVxJqOdpme+DUTLZV+tAQ+75OTslVecuV
an/qlsjirEIoEgjkyDipLYApVieGbwonUYsRULzmwKfpOyH6d8HeilsFohIkFMsP
263J0kzESwPd5+gpcTWEBMegZSijHsFoiNf/BaSsCPn/8KPLoI1xtZMK9Rj38t+K
YVr4L4nu/XpvF3afQISNnLpmERq88y+fXI/QSn8egKcMcmbFsl/fxYNWT4s04nMn
qcjarmAsjxmeU/NrtsCML/vkNc8xGn5knOMOQrITiIPwXKUXvb7VmQH4zOjbLvqA
TnDuiM9SMI3egAJsS83UTt4JeXTojN7Sax+p+a+8IQN2rqyvYTA0LTWAV/oTIt3E
fPAhFzd+mwP6bZjwhaXmVbcYHbLNSOp7iyFlYTkdV22M5lnD/M6PticP13L5LrjW
uSZOhUHUH+PBrjl71Rztc1Z+JTDoqwYUhAYZ4xCBwkY9sVqSV7xEb1PMK3aiaUHj
WStMsJ5i958YKGn6d/fWKop+JoUpu/bQs1IGgXNdSEDCStGygasLfd86of6kBcpZ
P1FazWJnz4E22Cuk7kzFGQUGPsLnpNWVjtQIXXdAV2zVnBi87ZrTZEdCIFu+uwle
gCvbonmDbwwc/1arvAxMiDfisZWH4nRhe94Wn5tE12ab0TPmyEJX97wbXreZHaso
7osHxUMLiSJYBcrztOtR/s1UnsRIZpRC/dPIlNhJ/mpN1BcpvYnwMWoTrk38HQfG
RPbL/DvpMPqvpFhlgo2FkdS5ZrfH4WKJCERre9/IwQSaxpooo/g3exAnxJ666xTp
dsAPqGGySmDaEVsarZrnMjtbB371DSh7ckqgfom53ZX04h3708TyhR8eBil+iT2l
AEE/i9vrpGDzkASluMBNleE+e2eMUStdtbicHkQHq1ZvZQO/TND41cWcFdYLv4ag
PblzjsPz7XtvUbUq3RcLrryOyDuXYqeBbPs4ZMiny9fcR5FxBekwvWK2FOHr/BgP
z5zTGJXB6x2tdUVav7VlumFmfEhhGAf9EogT6prmCsJDn86cn4XKD6ZbA1oo7H+K
4Jujri6W6HyqOjv5dwK+mJEA2Dhdzdl9j7i7dh7bI6dGJp0jST97O5GT42rCxODd
5yUUOBWSTUUTRcWXAwozIbNRZH8P7zPtpgScPVMffOF1kH+rOGYq8QPi6DAoGLp8
Q5J+8UM73RzjVquAnGqHq2BrTxjjUQklLTEntK/tebkuk53jtXm1B4BZDk+S6XRN
iM56ege+sls4g5PO5asy4CjHzVOJkw70qwYfPddSredAN941vur8fM4jIQI5B0i4
1b1+GDtn3HINmmhGgHpixVOWpdvsDvZEW/oMw6qvZZBWvuHLZsKFWM7m3MABrbgR
WkkHxaDdvyZB7bAnep2EYukRI9M0XLQkiLS3BAHnnzNhtCOhlAx5bGzIc0DNTTd0
W1GshjOTy45NsvPzXsq/ZdjDpz06hBwRFaRJPZVRMhqS1DF20PlLj3tSKpordpNM
3kQwvOKzpF4ZHIT0jpqw3/xMa8kCSIajd2Qw+/DRs3GXRJfAxcpXmHtwr1++7mKe
031xAFAFQ216fePr0txwtFC8/QbiuFetQ3+l9itV7DTQgfeJIeqm3Qi3Wiv8jiPJ
c0R5Lx9ST4LSWxvT+1AKgYaVLkPMjQGhk7LTsxph8CR/L9aeMse2Hk8Tl+gXMKZX
z0apSvzl6Ioep5hvm3UrvTl7iHc5yh72gfKbKxi0RmHemwQHM133Vg+Oj1DqCy89
t+MEKCLbdQuVePlkk5uy2eP8N9g6K/N4xIrXRypJVm4hAP5EnWlwJx9moyI5wfq4
Rz9rK/LYWqUnQh6AcyLKKimvQN2dy4hKbYpikinGilFHwTH9Sf8sHb0LSsmDy1ka
SmRUsJYFtGXGBIKvNhLxie0c/LCiKgFbSacp5qvAkakM0TvbZ9nMUPrEtvB2U5kN
hAzwU46bPWN3Tc03lvMbdOrWNbXYF6kzY3L0uNBu075LxKox7rxv+d3xgrBLHvzS
Kie/JI1FNQd67yc0gZmO8Y3d4tRAsd5GIGHGSpfpqFhm9ZLwFhkPUEI2fadLU2eK
hhyIcm/NM3IEFbGXkJFGzP6FCIgC7a4ojMQ4f2DAdUTgCNjIS+umKOHBiHHSeTCO
/ka5chZ6tR6WmleJtW3rUopsCZmJ5ODuJIbY1B/sTp6TBt23AMcNUyboB7YlGwb+
VeWzEvXOfgC6b9/pOy1NjC8+m3/EzSleXTvocpRs6CgIomJ1tbeuYZQ5HQ4AdkPt
N9GZqkxoM+eNbYzV47jtEQv2MoOdDCb8bhrBJXERa1RSFdQ9hsSmekwEbkJNWZ/I
jKRkcZn0oM5Gx0hqBebRD99UxJc4jNtLXN6iLHrkPZbQX2lnhdYkarSVI3CfskxO
gMbOMCyeIp7fVlAbdto+xWtqL5GFxV1rrBLRMzNMuv9N4wB7Rj39QPmKuuXDc2wH
PmaM2W7b8PGFi8Xv6kerEElElYF8gyWwaX4yA0kETsSqHV2di2OkJLZXRRsCit1S
cuSVej2Uqf55y86MLV86roUMyhDPPD8TcI/+1aKrrDQS/pLpjfACZ/j7hsDs8VBs
LjdMftQuZhDBsSHW/URtAI6QY9v+p8ygm4QcaC17lX1u858WDyyZW5teqcPzXIPG
9V9gb1m8tkUEYiCknTSw1Y0XQOZVv9OJEOcSPgeBA4XerzCpfDfS9ZnCCza0W3Ud
ZiBHm/VTfBEYPbD9Laio7uToxMRtf9492OID2gUG4MbneIAHjX4Lx9ee3xY5SsPD
8XehTx2J2reDbdGbo3Fo2vLzZRUBjg8R77GpyoGApOrtgfaCQDUMGGWqZrzPSRU9
iuJDr0jneXaJrMwf9fwb03ak3oZt96NnvR5vLwrNKs5SygGeoidLwEaBfxGgwTqV
rgVNWUvpiCuNBx32qdYKHTFywx38b3SkMm2IqqxJDcHAV9TuWiYP3saTijYr0XLT
Ey6h213JC/kl9Z7FoORaQ+A/a1x+q9rMYay4gf5i7/DLju092ZlrdyqoV3vIzgNV
GtosRdr56byAO5mZHBSL45H773RUOgfoyIZLNQCOv7AUcVuHqWQsojCbI86L1lr9
BaavVpk8C5Ry3yrPmMErAz/Pb8u4136hfp/ENiJN3Um1Gqygk85V/IFRzsyDn5tz
fGhMw5JJa3hfktcPc3wH/EQtJrmL4xsu+EmLsmFTwFHMzfW8Yc2IEjc8vzRurTnM
upUj/VxcxbhJYRvaSGaE+FmcS7WhMtPxlQdjhgL1iX0jwVxdLZCC79/6pLXq5H5K
M7LGNUwfJ2hD2lnJ+VqWSdkp6VJFSKwIRqW9NbJty+ZJpMR3iUnnvxuPXkLzYbl/
SP/p8gXwZI2XSA8k8QCU1C6UvdN6Jt6voet+rGTRJeH9k5LomVIt39TUZD46Gt53
DD5ym63n73xQsxUWf94GPwLJsCPeUKMCPQDNL50qFHdp72B/ijr0k5S4k857+zay
WMV9OmV5gll4ZJiUKtXH3Rgr71J0/vTdfbaxeXEn2O9MX3L36QjajIu12TEFnFDV
2pBOLqsmSry3La0l446n++GCYPp0n3szI1o2WyzI3Hs4sGf0UNhveXYxL4tiHg7i
qgYA1dHFGF+MLAMTJM3cOMsx9h7Z8KWGeNSXXBnnBpjNv4nnuTL32DWFE0Z8I0yA
Go9lMG0SjFE5EhygpLwKmZHUvw6Vewa5wfPTMZ2yuzu/BIMvKldXysKFyF1g/Jde
vuaANfS06csoXJBw23/V1DeIG0bjDVXjI3yeIsQUZjE6h9f8fHMuP2xZHSWpOguo
k9DWHhDTAGZAwwRj8OuDF3yFZQD7EQXaX6DQX9IfsGVKlGW3OEVgaSuKk42WxoWM
UitiYY1kEN8SPvkigriLFFP7jQNfsvvi/opKDGuZ2CVKVygdHYQhRe/gvgENdnGi
zZTxzEN8oTi45bzeWasLdbC0B6o4JFDkeSy8uiqDaIovwRoaLROItQG4SYBh10ku
fF7RpDX9O+QTKu4x6pxf/2gEmhtW9fwetqGOtIdeQQIkpMhq8KiV9KzwMnKsPT/h
MTKY9zVtu3R82o9D/HbPuWvewd5qT0TLEviEC++3bNYlmXEGD6l3jUmp3JQaO1Er
Sh70rItpk2wjfJF1kj3uVepe7cRzShWQjTQgsa66UYw8dUF0sFFeyGY5f6kzYVD1
bRLbjN/x+GoYkUdaPPMoFSHH9iIN3h9JlmvfwsBWlZLpzKxZV7oKvqfGmXi++PVU
N093Koz1jSP5HMpflCFAA5FDfidJ3zhDgNDZ1ALrKWUDVH4H/ZCAkW8PPdr3rhZb
WW4yyQ438DbPwdaNKgY0agLC8xDviHB0oS4yhZk92mPiY4jDnUf3reK50sN32DB0
NPX4umz3F4gpl3LKyE6TTz8liE2ph2kesTdfH2i1Y15HbjBWG/ZJ+uYw5gkzGMm6
QF0H9HpqnMCwkrmC6qZOMj/3ow3PQkn4loutSanghnFX2k2D/Bcs977bAK55JdNH
UQ6UWDLGWvZcN45y1S+W4R/hhDvFgitoLNIB5C/z0RROHa9+ptQxtZB/JSEAhyVv
MwexLMcLz9Lfzlky16iAfE+mvVmYWWDnJRDRkuGz4yr2HmH62gancDZndSVB/T2O
jrgxgBO1DmpKfqHaZqStEoFQIrxGUq6y3wgibeUZKidcO5FgZ2S2X4z/8LfRWu/i
yxg+NvV8liq7fhPurk987slPdo1ejrCeuXkFQQOEsJQpNIhusrZoxwmyIFGoQhfM
tCrMvN3NPupbfJGQsE9HJTZtDXI8TVYrY6d1GSKPCbqFQk24or4wO76K4qssRWd3
URjTSTajRdLE9quZZUhizO48gvOTf4SF1YXcagvZU6UH5sWvOQ4GCyvwIXq1IT1L
/ekbXU9+b0pd9nejifso4neESDlAwQWRCeKxRDWv06iDyovUKe1nZOWAqUMrbC3b
VFFsiMrvgHWTCbddc7nw/9pL+1fbt2wZAice5oa0DururmurIZEKyfXlrp7ro8tj
qGQsSW6nyJUc5vOl7hbtQXrqq/2fORpfYxcjjGp6mK/gS+zJ4wmKuBak9wnozn+c
oLpSuje9t6+mPvd9rXrkOxZdTc0YK1lD+VQFn5NAyY7LhuAiS7u2Y99vh4g0rREw
lSvrTtHnZATJKYuvd8rCpaSfLOmkibOe7dkTJqWid7yoFreYzSb9IiEpyS7Etd2O
y51VoCCWab/pB61PHxSDr49T2HxAHvuzs3FZmdfhvy+Q3CII0EFtFfKYBXDqGqL4
yEUOXqNKzuuky6J8+byGZCJy3qTwcqQM0Ea+hSDRly6mRrA+CfgN95j5zc/070dt
NK0FqqZ9WEuflOwa4SPtGyv1x1bZRRm5GFv9dD3XAEqKcJgX5aHUjPYs2j4Z1EO5
aua3PMc/2/GsBbK/R7AXmuGdr4KnHDGdeKMd/jTKEeGRvIK/I1Xpzin3lV5lUbTg
KaacR7P+aGHBMTaFIYYOfCFKjWqyw0B06Ipo3f9sE1uM2VbX1KuGjNGoOQuMQ3Fu
2VOfj1WOmxxV8oQ7cnojn7Id9Z199/75ra9tPZ7VFOMeYVosdKFKZbi91RM1rNr4
rkicTN6iQUbU7jcEb45MOiceGVN8OSluwRYGmiz/bxLl6IUKfFp6RtgwV/Edw+MP
IHVHWA9w+dKdoiAnhEi+4GR05HpRT9qD+JmRLFEkj6pLz29GCXsPruw+CMe4aBEw
UqmklGvwWhcAhVIHuZZIxQOteIcGSTJrptbAVqwFOfGt3y/e8lMvSY0nkzufZIYx
tpypfBEAIhMdrVe4rSg5alLW4omt2iqxkqONzVMerf6GrzxYAuMlIKGxaPAedMVY
PxezfgHHisPYpEh14ahz1ED2YkByIgaHAja79YEiO2ShgQeKrufPNfqJ3NThAzLO
7GqUXWesvzBQOd0wx6qAsfJsy/tkblkooaBrCp33dMZXiVCyQ1360Hz1gl5e7eNo
YdOQf2XqM7IUICD3tOUnJsiTgOl6yN4xK+A+hU/pMu+VP+nR4SkwhglY8jujfq0D
8cea+LaeZUE2deoTQtCxeRIFvRPyksrrq0j70k7R8V/N/eklTvymew15ozFDpjRy
Tjta7++KmTHQ9pk0YjvgYUzZ+aGd/AjgXGzYvw/RCl/yLv+EoF/geRd8uXSgzo7S
C6F65Zn0Vgr/N4Tj/MurPXgNGoVtGJQT5pPDXGPeAAxybwPKqHVKpAuo4f8xZZ0i
936mRNKoqokJWznMjJNF46BGWyct0fxJZcSllG/Od1Wya/AIC90lVKKGJkgrXizm
Kp7DmG7A6j0Jhw50y1IbNx8qp/F2c9sdfY5HGdwBVB163l21GOzXvF+qpdmgRHX4
3zi2TVBuxEEtx4PIMb3V7eTvYc5PWAkfSh01fASXbxL3Q4AzqYTPRddAO2lJw9Y8
OnN5rTY+kPoxu++JRjv2a/2d+48IO7DMMCFV/FaA1FOErXfxBD4FYkNQNxA6p+tn
CnbhJj0HEhuxnu7/nC5TfFpyFwtYrXbB708341OI8EdNWllvcgIf8YywXff7Pdt5
JiknTXNpVxOoHRdem7dNvhO4h/Tcf/IA4LDzBfSLWisyfFus44TM/F59NfABOTLH
qa4iEMpGYX/5DIGCF/r33+puG2XqwebZ+91q/YpunFnQHpPdYlMOEqg54fhGpJWM
aBIwomjVNLx0FHA6vYmjGtdUXXJDLdIM5zuE3O9ZCoZHY0l9MYeMWaWJGLDYAnuu
i9YajNrExcVGu/Pkhgz9Dsis2I6FGn5vlR9DOluU/7t4XgajG4GLmaCpPowmHDu/
cj8Yl5vLQxvJQCT3AaQRfoNXptuxanQiOm2EbL/LGCsZAoXBWuo2crS8DScSHk15
kbL60WD8fDgCkpJyon34IY1d7uE9zX/ggn8UpU0jLMp7/q8xw06T10JgNZlB6j67
kOoKYyibaiPP7qP6vyXYf44YR8M0w66oPuFZlztsr1YRkRqMBl+nTHBdi8raKMDd
fLTVrTQQEz3EHzoib1Wdg6WcUUw9olwB+tCTvJZzVDITuLxUs2jWVZQqotiQmGxL
GLMmuZ9M0ZX772Z6sfkNquGxlV3wkbggFPsNeh0lnXMRvia5vg5QuUPigB/7whUg
/GiZ86CRxPEvgZPjGqfclPAL8VwcAlfMlXFlO/PMLO1o2yT/uubqGP6Fi61bFoBj
Qg6JhsEAqdXJW3bWcvkEa9KxvIm7oZhADbMu9N2S+wF9qxUh2a7nfdM7GyrnNPdi
3cFFTFY8rWUqlFjtNYW6UfxcwVsJAAwxlUmScICRXhIDAEVItaLVYDsh0KCUKtCq
vh5AOrFWK3As8unG1rRrsxedL4XO2yQwkSP16tLil5rBgcC4uGqhWoLMD3zFuHPJ
QCjjJ2NfaTWFIkpHLDrnOq0g2ew9T3p76YnK2NX8TTJQRrgdTwHYg7ZQ+uZVDJh3
8OwiJ/b6BTWcG215d/sOAleZHGCCkjHPeN73bYFqdf6vXkOo5cyjFNnvJNrabW69
VnYlBa/bC0+rVGiUiOVdsLS1dNyqXwlu3ATqi2WeVBgTOcGAsKg6AqSk8OMptDkH
p5Lj/cLH4tqvdfyjQ6Eide7rqae/vfA/9xD5F98tCyOk6cmfCYp4mNXY9Qv6r40z
YlIAN/5K9g7vlK4Gav9NK3pdZbu2henalJjPgXyYf5SvYxoy+XmPiHkq9koVmkDv
DspTA1zA9u7xAC7aQSXMQwenXYvFm9RjyBaB703KeSKjyLDp2jLslQeVOItCZ+Vd
yumZeild213lM7UujFRFnVEx892hypt8GJdevCnszkp9BMSmEsp2zEYFA6ZkFeWA
1hhDf48LuO9BI7L4p7C5IX3td1z53noedVUH8Rh69U0xWgiWgIhxhOdrI3nNWIWm
ARz9GWYwLE3gh3wFz+sJOj+ukHfDR0inZGuBprr2Lc2Av59zlvHHNFs5YeQrWPiK
UZHURLcc8MKZUprzruC40HaTDFNFl+l3E7RFXa+WOeAzNP7QoJXh8IfWB4jjvO34
ykEzdRcik4/f4mzm9QSU6lQtGNUIWVixqmRoN0H+AgL0N7jqFDormDU6UBWjR7H4
HbE7Emmb2uM3ZyNSqffKFY5gJJNVnlcAig6ktehtlkUkoSNtvMOL8EJIUGRe7KNE
XDwS/vC7W3hSg/M7MkluZ0RgrioEUaQOSxqvoGjz+/j0KRbTCMujHr+/u+pkeFHM
eYPVUC4im/k/m9RS+f1KsLh+b8PjrQk5LGI+zrfzVnLw2Krau9zj7JUmMkVbk46l
Pp5EptKEbqnlzZXf6ezihcmSY10aKEzRNcT629a1JWev48UT8wtKYe+XRRfnLcfL
1YcvYihtWvzIFSjvLmTA8f8sooTl8TJU9xtl7/NUNETvXOdBjrj8MeW4qpPNf4go
pXWhz+GBzUe0ODThZ7oqf6Rk7B6+iMjr3O1wOesIwioqzNqUOTUR7ZCH7JlgQidT
37tIf9WXBxIBtyBLecjr24qT91/vFO6URtZ02efOJQ/mJZHHeB+T7UmyWK1Je+tI
8YRJy+Wq1+fUs/O1UeGsJ5AkkYPdf2wwx+bvz4jQ0oDeOLGQvjPOWB3JGlR3GJlv
iTH65wpkwWzCjDu6iX3akwqQGFCzvYO/kLX+BoXXI3D9BnU7YujXdAiBOTPlf5fe
e17WfLCyJZ8B00M8QLl/de0Xrw2rp/mWqkuWkF3cCO1Jw89UXk+SO4cVnqu9LVi4
Oc+XvkmH7KORcn6AO7riRDz6p8Qjyzbu+LzfHSZZ3ibPkb2T/AX7mDRs7XRnMuyi
7UehFz0w9MuXMJwZigec2tZD+R0R9JKRA6VMQnxxG/aMkqw834ylp9qEdB+eBFfD
Qa2KGhybP4huUg4hHxH056eM+dB6HCPeDlgg2BhAoM4ZGL3n2u01xd7BjE2TkiVc
RggLFTmY6bKfy8cv9FQ3rBHD1GS3lJYK4RcOhmirfZERrjdLAvyex5tNrwJGAuTC
0KS3AMOeMRK+6YJFJTOceKl0pntCIHkR9dTBv5KeGln0UbrKb23MlANDtag0Kk88
eeEcGMP2IR10xIyfarq/KLlffQSQgp7sN9U/w4LXIKsppHIuVkOxLs1rBG7QTevL
YNYfkG7wbmQwPYmslycQUz3UFEgh5gTv06dlfld2Di+SBmNQzpC2xVeV+zycpGhS
wnejX8/RbOPn1raiS5Qpte1glSPRqPKVmstTCY7OL1tnGUemlWv4t+do2djzwZht
CAJJlDQzQx0+QWdD1oP7V6TlgfsHtGxS6l9lNG8YZFEnHmOHSdVi6C8pMZf+AfWw
b4MkO5uWl2LAteZMlyLlfrHWW+1d8bohSRHgmGz0whvR0FwK+So08r7m+jR5nhpF
mSDjgj3QDSIJ0Oo2aw7BxGTcOm2+b0eQ2MoNUe3Wz9pLZhn2h8ZxSVYv4tTP+Ft3
s3xNV5GZibWhU3oNcOEuAnJ6gBTbkwGUybOr8aCsMqj7udXnPbbV/RNq50vd6Ix1
TqEOk7o6/2JGKQazR3GEG/SqAuwA2rR45vLdGL9ELSTLuvF092haPm/W7733M6fd
y8x6Oq+YBkThC7Wp8WNyty7fVUw4+UW5HHOc94Y9auUKZlVbSqAKCAuVygQ8cDil
mBeqo9Eefj/uG4ZSOL+DMcsVTaeJMSV/zLTYyESJByEfacD5F2WyHkhdTPVD9D1U
+ahAXLSjW2zhGFnUic0p6l5o92Z2GySEyTtni/rsJshadB9Y8bm85Ipb4hVSmWeJ
UQOgbMDul1uTzpoTUalpV47/GC7eoJbxBCSZW+svWXm8xS8u7qmly0J+Io9cpeAI
k81NXRxQhzjzFxfBqRZJoCkdeltKdc9yJiJSC9to2HaBBu82NH9TGD4MJwb8lNh/
9Ovowwl5HYyWLrXFI5jmJIg2ZWWHopsGf+ZalEct5o/fMqzn1r7kXA1J1oinGL81
jaABl1/925cKx4FOmFPagGOhI2uc0CAwut2YyeSBld1VfBF14R9j6ep6PAdRDEJF
4y09lqsfADofHHL85dd90R1LUlpg4GNzAwTEhX0tJIyqMVrsvTnIHUrVIBZP5+co
j08BfoKcNY0t6qM7vHcuzkAZNUltV3DqnW03/TFHKd2VjKWeOzIItZLQy3tAI8aa
c3l9OtTHry6/tivjuY8uVTGffO2SUGMvSKGXxBWlEsMvzZRn573GY7UuUMiiL0It
CSnhpxS7FlIcOhMDM/IjxeEKuhL/QJUDDWl3ywG+9DosAeJPwP8OR1ny3SpJBihA
Z60HpLRZEWuNxEx+VwDSkkdDR6Kbw12XdnG7F/lMxV2PDIEbFsVMYDoLTxj+5HOS
89ssaNWa2x7VowIrRQajeeaweogZC3EwrvwopcAk5QnWLOgn/aYcBzfWzJiZGzHT
90BR35K7Duyb/Lka1NPw9gQelKU1rLTNfijo7NIMNs3dDAmtoTDCExAjoBGiqdb0
XbK5+Hr/MEDrV9qujrSdogcBiCFTCa0ZTkPaZfla8BrTb2D/JVQn7/SdhfTdtnJv
nRTOJlg/378YjpzLO14MoiB7Z7E4rDEPOsEEjhTVCC/7gO9fOf2Y91xigLJODKYT
K3sdZN1H2b9uZE9bMUTHcTrYdfnja3QBrqbZEs8lyZg91rbmwfZbOQOWl/YeOFr6
IZ5na/3OMO1pkKgKWjL7dUc9WwBabGGkk0nwVkoIwonqWTanhh34U8gEFvWJe+6O
iG8BPDYETRiUXJlhUM/aOOU0muNpXVILf3GM6BiPJPPattGcuQZ5QvxYmCIc+vzU
S/F3ijokcjqWghAqV4FeBxwfH6743Ll2kbbNKg9u4aNFGZOH8HOpVzFbR9NvrFDP
9+Ml2rRRwYUuD2vQSc3WCPB9e/L9nzpq606ENOOuyJMipvPynXIJZ0RRIbYOYv+O
vfO/y9xkC8hNUwSdB1rA4J2HDxhgTfs7CDI6ogxgX2nCuzKJxrhA+evZr6hcLjj1
uqp2OfKsbupC9ENeg8rAxiGij6LbaDm+PnTvbGx0U/EFW1CXWpHkd/mNjUhjwX4o
wbLpnqY0T3fQthBElATGgJYgE1uYInk5XB2s8o2pkz5GyQ9pisgL7ilrE/injDKE
TQ5Ea+MV9hk9eWxd9gYhX5jTb2Vo7TtLmd+rfhVrkuwoA2j2FGqRWlWZec8HXQXX
nFvVKeO5ZLxASDxcCb/GAsnJrp+wHq9IjhQKiO/f4zdQH2SVLPFvEomd0pXFRZ2W
UmrROSFDYPKVDJnNcQ5Pxusg6gkcdwysq9OhiPXH+/w4LlrXceSm+qRTXYcfU7xM
z+qI0R+pTh4HFw2QHx6BlREAO+b1ADfWMGHZQFahHaikh4C3vRX49ub7ibDl0NR+
kvL9xZks0D46pryEy3+WSpANLYMDFjePzrhIWs4bfnqpncZ1Xwf0FvnNk5tFaRHD
d2QeTmwadFNkcEu4rzGsobq6ELrCmHELdk7s72Hwgr8qS2t+nHbUfcRJsLo3vYpm
3W+Dewle0b1mEfLVv+8wHRt93qiquBo7dcc2Ws+iESDWTij43mv3vW9ewC0rZhSh
cDxtFwyCcifiFOj/RCJV8yy1D9suTyv+ke6tPrUqN7PT0hW+54tZX44LfaRe2qU0
pS5DzJiQjgnnOvRdOPSvImzOtd2EPPSfxIjWNrWlvkR8+NidXfnoYrIxIwuP3i7p
sf2zrSPvNPogWM9FemTEcc/8V1Fkg0tHX6uQuj1GxzF8uakq7WSvnbpjYlhHGPdg
cK/pjoa07EQFVa3sai4oOVNgWIMWJP36zx/zM7axGXlHjcti1QkOMMXoMhBTMc2h
3satav0+AFIKsNce2oA/bEu5xQi4xld2p0rVVwr65YnGCYVJH7Hi1MxIW/loWZUv
zqal30uLUmKzx3ktZe2VPjM0gNHn2ArzbsqpIcQXXLMwOBREjorpj9Wp0S7BvJ1f
EOO3vrpwM47rcC0TNGOGOkiA33WOjh0eewFSy2rDfLB06C5drSXd6UtlLj3bzTLu
q7TxFFnjQiH2FwDWhvt90XJ6i4jom71Sfin9whOMpRUrvnjTNq//Z3NBdXqsSM6O
0J4sNxzEuswDSsYxGT2UKm6Bj4KQgOmCKs3b9ktiWziljgT2qC80VKOBCUJAQgLe
EyPY+OCASfUSZ/3wkCiwXB/dXNt2Tq/IIogeCfdLgoSOFZ7L7gOUV4CrfizjSXCb
tBu3XG8h0SuAsAWPVio6XvhXlyFiuJtAwAzzxSII0giy3bPI450pyN1XHP3XQclU
IzUZ3rSiPbpeSII4/G66u5l/Ac+fyaGpl7fGca3ZyWnZU1sROt8aZt1foIjFN1qW
FA8ENUrrz/WkiupichqgcpYzKHCjNP51fHOroxLSU1UAP+GWTHtoD2YlgFVRPzrA
mSrtozk0NOU7feqKSz2aCTtPd/tZ4Iwxx/Gw2iyrlX7mRfk8FVz/QgZD6ByYGpn3
zD/KuwBh7oh0E0wSq/7j45Uqbr9W+03PZQCpQ2NP8MVbxDHxe1nm7SUPmZZOKTsb
r7+3/ueRH+j+EE6Pl9Hl8egaVkQ8qkrDi/lly+E8w+CxJ7eYHyIbjHLSlXZWPpcm
5ZnlDHO9rhcrGyDHZ1IDy/lv3KuEBC7+CrA/tqZineFfi1ncNyZm98FQUWKktVIF
LCl8NYDSdwm3oKg6Sj86h5+jrTeAOqirKdKr5Vlz6J6sPQN9kJehWpFLTvXz+QLr
TOfufJnPMnI6Skv8WctrCQgNiwwXDGq3MiUdbQnAdzh6Lb2rnmWY+xSLYmxWXTn9
7ldGK4VHFPsgjFzTFAlHbH9BK9aznPTddcq3Z2f1YVaUinvHMagdWNo3U9Z5Cu/D
UMQJF0MbAzWuJW6ecB9J+7d1PERaNpHaCJmGM6DFI2MuNB7AxcAGviTm0T2kUfAO
ReLvRL6iW1b1W34+TSx2OAa5WJ9Viec2E7rLUhIDBugayzOriBfMJ3jLfTTozbew
gHsFzPymHlw5sR53PH5LxnRcuUqxNv7oYNwA60p4n493g35HWlxUMSBud47rENkR
Dd3UiwqYpaejIjYiVIglEYaZTlCCufGpMGktVDoAkyruojwQtddAleu0Irkan7Wc
0qgH/fw3cVs/a4OFQax7ueDU3nn9LAhNjMqG8XhHtwh6ZTT0J8KXPj5XNxPlvqqg
bIFRVt8+UF0HI3jghfoqg6yaXmRW/mmeIq+swIqD5g/gwuN3w6lPVOTIl9ylywTE
Nqojm2q0NKG7ZT6qABj26ADhr0JqqlwwK2QWhpX5D3CvzQkXu/Xt7ONfeTqIajdH
50+Pwr9Q09sCNrCw5Fzc8ZY0NdlnC1fugBgqgGo9/wFZNREo0ugivJ+4A+htL1xO
SIvYroKFUD3jiBTK4o/H7whVmvUQOLTvmLpC60Op+IyjByo1njFoEYxUPJG/S36u
UIRmycsT0PkS69nafBREmzPZ88FKBOPK0ZyFMXndD5jXKOIK3DtqS342NJUmSRz5
QQne8D6iNr8KoYiGnY1fAjQ1mKTyNwbzSHue6LKW4uG58cdP0MGonasBmbs9mxLp
3dxL/kKEX3haIeQ1T9S20Hx1mrR5OTLIlUJitdS7q967cJUD1L13Tb0FzViq+sxg
Pv3Px1+K+Wk66I8iLV+adHFdCiIwzRnII75ADhYMxJz+5lP6CGJFMULPTYezGKnr
uMWg4ZCI6HVFlApy/VrhI3WuSirTcmaWjUNN9MpULulMDd6D3wpriW7cgU4RmLyJ
x9aGJZjhvAR2Kz9CNuD65Gb/IWCQFsBvjIXUgPWIR8e5ySCK3/VBizX/GbhrMbDh
zU4jiJO7mBK021L3HogzaxydFUywNRyybMvpmwzM5oW4kvei8RKiyfq2L2rQSGOw
TviUDDugnh4mNtw6j5lMP3ph4WCorAsdq6bQtVEbL9VT2qMbikNQQA4EzYSsSAeS
6dxZBEIG1tQyuaHx9FWg5OlqgMyDgAl8gA1/QrmS116WdBJouWVLzDc/EnIKK9OM
N/GKCPb1gq8ta+7Dl34UgChZkSGOo9HuijB9EMdQapozdsZo+xr3WBYxsBvw6yuo
IxYyhxuM5lhJqYQz8FBiQrITSn+tX7+q10sBulnhN5UvTuKyyX2HwnTEWyOmsj76
68UCuEFZf5PLhhoQAlA5pC5TiDIKF43uWDlj5vY1Qb4+yjF0ehrqZsy8GYEH0EuT
/xOLtMwF9ny8/hfDFcQ2NRbHtr6uJCB6se2tyMFlzTDRyMpnPyyHlYj70H+EByHK
ladp0GaGz9cx5K9sfO6Xq5GQA2res7nQIi7dSBorT3VaHgpFtXwV2VzOt0WtpWsU
/lRUHVRwweVVii952gnKKOqTExfz0dG4ulxWMsnFHI0nfdlimP2pzHcK7U3X2a06
D9DvCyuqyRJNc//AE00V2Quu+1C/jd2IcSfSdgohUIPK5CFxhdkgQ0rl5nHrUXJH
7ghqR27p8lqDhiJMtYs4omhViIdQTy0jbVeEvgsMAiYb1ecUxCMzIgO6yVyR1Ube
wU9Hrs/7CbWQsFHmjEAHDm38WVQTywLY16NA0L1s8RLe2FXxo5bT7ZqsIqqZdyAt
dAdFzcXZlcoz+nG7/73nQLUnHfipnV/k43vMoszkcj81iIuF5Rcldjf3E22TBKzW
dSopS0wdWC3huLOhMg3RPNluJEhLXe9hb4G7kXLg7M11R8CofMVPGQC9lSzJ3f6q
ic/E5IAqA2Gr7UXyutkMzfkrYZHZAkvwn2UdFpIm4rOxhSbvRWxilxCNdGjIM9/0
mauktpCY9KOT3KRbbKC7MWFbiio7VkHYXhJ8x0HnxK6SqXelWRGq5Hms7NR7Fqw2
qlG6N9cTee6CMWFHYUG3BMCPRFWvMyjj5UIHSuMz4EoWfHUDAyVP4S3cGlABxbF+
8lUCAmu6oPd50qj/gKqs7HW/Ql6TuPLa7rXJeWT/TROvSSQ95tCXQQ15+87CTeKo
BjIODbmXAJCdhjrBwC3CT2kDSU3AucwXzIok9NPosg8TtBPWkHVEmIBkNsYcmx2Q
K1mP5BUI6YVauKZMliutcAk8tM1EGv+S7OTrcVilrvaxAnfTu+NF3lcKTkddu2+w
UdGI1ETyduzrVgqYlu8PM8JNgOMbsxEY/hDc2lI/5SFY2eBrYW7h10F3qZID/nEX
4EPyPVdElpE+tVU0GXT/QOHcUR5LpFHopQgjMEqCidhun7epGaYx/EJFirZ5OEGj
3ETDX0B/8fnMMKK2JzqnS/19VNnMa6+uAfU4o6AC+civjktRsuc2dgiqMI5V9hmM
MsFB/ie4M+UFhh4TXoWOmhBl0SViX1q+JtroqNyeevr10pWwCJ7M2O+tK4mne36g
dOGDU3acxbGRqoencWMmq34gf56Ab+tPYrqeXSzBMaBqfnH1r6YHLjzFfmsl6nOS
MWvZCeTm/Xi7BLKm3IgmKmPdKxIeclRhi6BfErqz5/fuWOjclHoBpCXmAxSzsl72
wZfF7eETPJZElo7BgnwB4m6tRur8f+fxCuJ7AwrAZ00DKu3Iu/8/Mrp0ysZaooxA
EM0FSuJsu1LMwNqBQP7EW6qFM4ywPgk5v5MhYCdASZwID6vrPkLC+Cjvh8RcX+Gj
plRmc4MLIJNum4Is51QoAD/vvrCBBFJTV6EoOPPt7FiNGMu26ktA+UT/fRpIjtEH
pqFFMb6VR4tA363VzEVtPDFfJMfcqOtP8ZmSpbwo4HdxXAqZJEnpBJ0k2NlL40zC
apxD3CEgcDyXzMyK7YWpWZDO0TF4vIUnbpfkkBfwvpl7EU1JWkoQA1iFyIJxwO5E
tT3fXN87TH8/VujNb3C89RMMzdHs5wZzCRQoWVFAK5rIsv0RLxvhM9V6/A9PoAk1
2qrifM31rRSSl1sJ+0c7isC9G7pj9J1k7EPca4x5oTymmD9rYTPrpWLmMJlGVUdk
avbdYt0Vy0Ng120ScSnENKGfVFCibItWSyucyfT8H+Ps2km3a48g8/QOee5ViMcL
Trw9b2oOs+kOpr2lQHc4VK5jmUvBwec20hGqHprzs8XFMzWaqt/BC0vLQB8CTVna
OM4J3c3D9W+ElOrpMIVofj2Me3T4kp/DR4O7H9DISAQMaxA8Qb64kcNaACZftPJ1
9uA3qhDz/UPAW8dsaSEmmpfMHelmYfGeK+HHzeb7cXRoHGZ8NCLY7GHE+TrH0Lqf
5sm4u93iswHaCFwbfpf6AUQYqJxR+v0D7xaTumpiDvSjmNW3pKc9QY2QBPvVHDUg
Bggwi07OC++gmY1tyv2LlGDjbJ3ZUrcodxb6lSV1H4b2tipPWxMLiTBjNhB33V4R
qJwXcB3RjWeKOnvIADurP7F9lJjpr3ITHqqfd3zwPF/qcx4njqtBUv360GODwXIk
SLWK8grquUrcSDqzjW7IWbmuJ48j3nDZeh0nwgveOCs2ah/nh2vLPta30CKRhpv6
TXX7wDJFhiqVY6MSzYtngFE8QSshlyOWXHAIpEPeNHmtF2gztIL4yIfFBHVIn4rp
YhO3bSr0+A4wxNWXN/m+sQ+JAIYAJz2qDkBFyjajZwl9WUK0/5bL1hziqLQalFVJ
G7kBRRE9e9kTj+MJqRnIkkZYNUZ+/9LWwK18N4Og++dYBJmWYm2umNqYkh4QdJ+t
9lNt9YNjl/yGmGPvpeJE9FJ5n2LyHmaMNqEUHuKveg+1pTU6jFEicd9P1+LrbP3X
+/0DWJvSdqYujQLXD5z9LaDAOQSUaeC/nqrtrvlGjdlotFUZol/xzBg5MVufimJf
bUlVvatV7bL7NswpacItemdnuAG+vok+1UNHKP/EzVwiQb0BaDn9+pdQ+YgjBxjH
LkCZBwykeh5Njmk+1vgWBPx5p8ssefgBonV2BaY3bePruklyQC9cFUtWiOJn+CZT
AYA5BePaHFLDJid+ldiMgBcZbFlvjrb/4YseCR7jOlAhzPXQxNR8EmZb2aoEkbkV
NrSpwTdhxPXQHpMPdJiPL+OuNxh+5pcSnVj5MKNoq6+kaSvaYvCJ06QKGu2I4vMB
PB3NGQhm2zztrIlKPu3YzxIY851N6tqSgn78kXm/n9BTXGHApR5zz0oxn9A4HL61
9gifAt+uP7SL3r6ateWR3IS2LTpkJbpZtCPPjGGCJKx/55g1kdmWehJCwITB3CsQ
8u0Zly94b/ui8FLOsqYLuGFzToy5nImpBp+NqdvO9to8jXeMza9+MY9mlRoKnW97
TqIaViptSWFXEK840NKuQWr+hshW216LrnM64lK6/jg6kfKSsQ3vV5ZVLK0tZiB8
KTFEPlkZ6Q698YX5QAVh2k/BosfigNSCZp6rY9rOZTeFZnAzZZhmQB/1IsmTvfIu
evzZLf9ZqEG25349YmPjuTIelETbHYFZ9XhtQlOTsVkhLq1ziaLmzj31l6QwWw6k
pvB3tWwTvlokVnqBasMShsnSv8m00bdJkH52OLgEWQvQwNYwCapGo2jS5GybBiPl
QhzXxK4ebIFKarWQ9ewaOIUtVWhF+UIv5AN/qRVv/P3XBYDXBI9tiYLO/bfSYRZr
4tUJivkZ4sAfhN4hng8PgJmYqCQhoF3oFv6So50EQHA5DkvZyW/Fs1gy3DJursY0
rS8qsOlEZD3wfn41/RV498AssOfhQGIzfEl0wZ1fB6jN5ogPItod9grcdfZdhnHY
YEPUOT9ykh6Hth2MpOBeMEZC3py3VsESKM5V44+AySnh8cnxQewbYFGtAPCoZ0vc
42Mt8kH9QQCk+nXLuCQRyo4m3gnLQVkv6UsWzsTnDFaIkgQPdxHffF3TYnjjJwgg
6hipdejAImrglfzVpQ2Aur549YkR1XFCrGX6/uGyPId2mhcRaerRbYysu4Bzvy7y
7AFgkjDDiIIpJ5E3mMeSrgDEdqa/ttzjPSJO8rmieFiMPn7KDbYpZsRW72KVyUPs
H8vYvZnR8uc5c2mfy+4xnRezo6NGapGEw1zuYoUIPGfLIPvmBa1EY9OQFICCp8Xi
/NHITM3EEJvFRyJal47iAcjrXOtHaMDtiY+Eq00y+Xy5lIre1/BonESjpTD0B0vg
/Fa/bgWX88b3iTbx8NExqqNsUX2d+Pj79FBKf06yKscY4wl3I25P9+plJxOO9G3U
tdQYW9SK/iqfAhz4rhM/MmzmeHn4Hu/szuvgtvdlZhwNwT8MKLpWcwR2QcEKXtu4
CJVTYzqEte0Ogb3bAZEjmbNomHum2Zv52UEwh89GtGKu/YbboxZSvc3X3JNdgpjr
OYpHnDk8pqXAR8j7cA+XCkYmtB3WP5UrreROF8+X6luvG6Gy5yOAZo7svQuvSZIP
VAIIYwKyp3GOVgzU+pGEYJ6gIYtkq8sBDFJ4+gmoBkP/dKOnVsmLM7fL96wQVBcn
KtY3mA1u3tarDd7IvEF+LiYz9HCEyWDeenY7/gNLWCyFXvixH5hTtH3SKLiuBYPy
7osgTLM+1vVK2rDADe0mWN141qcSMot43cRK+MfBOSqtaJOVlGMCxg/vVA3bdL6m
fuKQNBihnl6u9b6kpSyB4da0IJsLOZEX2sTWVHlq3VUKWk6JNALo+3gBJ+H1Y7/6
qspu1WN35wgpttnI7oa9ASdUgN/2rxUDnrluN46sy0cLWD2vJ1HDBFGpBtyUTAIm
DzzxmbKKgPJGbqYYhP8J/Z9NAUavgvIECrdBhGIv5CCV3QTsUpBvOi1wSP9HqAJ+
90a5giHVDy0SyRpwkHIdi2pWsqh7NJKpgRnXSuQB+UDnhJ98jhGdO/umVB33YdH8
qTHd+nVrzLeB4zLHlPxVP/uZe9GOc/qzLqLB/guhqVOW/bmYM2plIGREV7ImHZEI
PGGWIEFf+QiSvC6Me8CbZsK7jTHMmnNPPBmKwFOlSh1kI06vipxqJNVdwnaNvOTc
1RVaCO7LwGxkZa1KR5r0+IAH2Mzjtvt1uUbZwu7F8fqVx6HFpXfOPZG68uMXWwxi
WpTQBiB1CMaKGs0BWZ4h06Yw7qmu52MMmbnyiGuPygjk+WYtdOSChZ2BiFTvG3eh
omqimXPmsHC3apeecJzbrF/itkATtr0voNKs5PaArH3IrWGcg53fuXKKDALQpjLd
tOqI4bI1DmhWCwnwDTLDU6gBxQvAwMYkEh4dQDEDomAbkpFgAuvWcauP8yT+eEeI
wzHzSox829IO5Mw61vKft5fR/Ojlb6wMPf6w60Gf9srezE9LKQu37SPd+3DbDl2I
6U9+GMUiSQu3Qk4kYoA0e3vV6PTt01RHsR+/7oUcH7qqV/O5oXYgLosvZdvM+lCh
243vFE8U1OmfO37JurqIqbDSY9VfGrtXRKM7/OZNSpk1v4a6j4178Tk/Hi4s5yuT
m3Om01iE9ss+E7ucD8t05LAVizOdGpr0vUWRQBeyXLsBmsMfKWpxU84PBhKy5NIL
MfZQ/f3+l+S732OIEyFinOeaET8XwBim7eDWFpOVHtGoMkDW7xKZ1Lpehf2zhSGA
IB/b12Ga3AHpbZqYiIB8ZLZ6yvIJpE8H7vy0ZqZx17YwAZpJ1NQ3v3RebsPcnglI
CgZOh95wkvp588jIn4f19/1xx1ZwOqaE+dliojRiokim5LwpQmyb7EA1HWwvBv4h
88S1QlFENUt7VmV7aI47hc7i2qLJbJfG3uImu3Pm38bK6FLenOm3OShB3X3gMkRu
UgiT+E0HHKrp1jwwQjG0HepKotvkcoSqQqotX3YT82/mKSy3b+2TZzecXzoQRDO5
m7rl6Y/A1j4X2geXOBXkkfM/x2CCJpu1A17Z2ZGEHdI3giZhFCEJqtxJScGyzbWU
eavVcYzFnYYkh53QfQSrKA5m1K14hcCbaI2MO7KU5t+sProx5FkET7MW8jqsqOaN
7EkE+iM/yhC0CJZmSH1Bk28ru/J80lQ7KqIz3L948Lc960w6j0mPaUkBEoqfVks5
a8CfWaiTF29WHAxYBZNo29eAvYxVI9cEn6h116tzl/oldMgrl+aAkWflrVQBbkEd
ZSDAiD2LVNQMhmwkjjeOTWteu33D7eJmjdpRmqPmvcrGYX8Z3grMpPt1o5gDtjhm
k3ggHEMQlJOmGZmrRQ7DXc0ewOQe0WWau9NQfxjeknKYs1VvwqL9vBUf1C7NBuTp
PflB17B22sUfpiC3wmUsLEpnYrsQNXailIUo9ENS127yxibDLRMq+MF2IRm0mUrg
6neZpHzJeZxRMJ5ZWkRN12YlKcR3REa+9uWWIZ9QggGb5W26Gthzog99Q6prtzVI
0iFTjUwzoS6ilFImLcrKtLtdm8fCQHjDx+9cKZ6j6DYS9vPvFiIbUtg1t0uCZcAO
KT59lApaCRUzGND+yIVjgQjCyNw3ttR0l2fs+HxUn3Z3NyF+ELun26CuTlRg3DV1
uCfoOZpdwkNkGWkPse6SHaHiAkORtEW7zYN1ukgP40rwnIdtwUQHBlhSayqtLF9H
QC4ptfyZWs82Y0X9/1J+7jl/NBGr+c1UEt3r1wp26r/YBclfqiKrdB/iyPCZDY1f
x4qf5NNnL/kkC6lLyj2LjOm1OOS9y5kbO0h1IOuPphHnHNkx7TQ9Sp5rn4drLl+W
MlE/G9y2q6xFoQZKDGKIPNGfvLUDQxhPcsF3UrTUNVxmofq2bJS9vDYC4pgXMBp6
68jcYGPDnZKw+eg6C9FfFrGDnpYVJEM5FEiq5e0YN5LYLhmjaQl5D2DEMBwyivFZ
GYeVf8KI/eNkrJnFM/fosiyKPfK1u1Ka/iXfDY7MYRMPZT86X+q1WNiPiOVErOPE
pSgdKkaQpJ0bUPFZpcDJNVuGNokZcuqGxLuATZPuS0spj8VpOEdPzLFvJe/w00FU
5UytPYcSQOwLp7Ygqwui3pVTTSaCDvSl9Dn7qiam5Wv4uR79ObpdTZpkPCmK+u15
tQYQoPBDvf5VRjFdNHxeciUMuLK7jrEHJC9v7FxcV5xveS655iWyhQ0qBT+EhMcH
qB4DcBTkZtIpiSaz+AYOszfqNUl49MEydzsiTVWf9uFbqCUE/5dYjNcTg9Nc9n0m
6Wzpg4ZbZM0Hv3eGPUX3EnAv2/OxAG/ROYxkVYG4Vjx+a/AemRiA2tAVB78tUR+v
GKC+prg2Gy3DnCcLsOXb2Xj1pUBBh7p6S14QWJi3OKqJSV94AxrYTuyFdMKQeBtF
a0Q1gwhxRxzgmYKGNiFYpGX/B2wgwGU+YvIrl6XOMytlbGDYx2dqlL5PnR/DR2dQ
2ws9HjUi7JYkVCKm8EovYbm0gVsYjzyUC7YxVPG5j3wSOkGgzE7TizECEhHMpLyv
/obdDbvoaSqWLEpWZEhmWP55dNw17fV/koc2av7+B96pSB9cUKopVR7auwzscH7A
teYlg1w5PBwM/n+ePEzKoovjNMw3b+PEF5BWptd6X49aeZ3QlD0NQ0iBPLNEhSvy
ExhqTcAiIeNvEKwr1hOWa9e11ZOq6Qc5suXpGqZsxKzv+FA69YQPWoy2qpiuourJ
0nyY0cD/sGJ4OVKLs7ctLqwp58ME3tAy9YW4fFhDOTR38ISDUu/mQNVtxb4enAZI
YebpVWzxf3Fgga2yAYDWugM8hwFg7JkdGuKxm33Gg2riHt4s2QO/+rBuKMp/TmWW
yGnO0O4QlCh8to8z/TTmmGn6M19NUJZvu7Hi5+ImPkZFGBIifUV5KV6bZm/sp/aV
OR7NWUfe2eRKfi9IA/DdOK2VUJJAcL7QqmVdr5YHZpksjqbEpbozvZnz07G3kyI6
+kSY74BbNHbqARmkAZMZvWQKMwfYO+ZZJLVyg0XbLYPfzM3qwzv+/2tv6v8nbkI8
evdH7J5fUnDqmS7IWXU7Z4JuTVEZLSKmS4RYse3bDnMZTZa+1WbaIh14fEOEHt7S
g/SH3RByaCfMb7rftZJkpz9h//sHVotInq7AD6OfqLAARxjBlobr5TIuQfDzBk3n
BIEydCW5Rbn6Sk1ze6bZD4N7ynM1eV9cDnxm2ErjUP9vFl0apSbBkTWLdtNjdQlq
WS/20LjKO6lQ1DAEj3DNZ1AUqkXLAJvuKrbYISNnnWYijrOdN1fAZO6odbwuJjYD
wp4zrllkn6leslyp2lVOHPVaA5f5adIC1xzr7Ka/KSii/4a3+COdrwkOopr9jRlo
PZyZCHAf3pKQsQzzj4+Tt/1jNhlYUsYCS65P7XZraE2S5YP26pQBwxQuk4PBnAOk
e5FTRW1Pf7XA4Fncw8PSw/b3irFUKIGsbxtG8mUH4d0t9E11dTldwg5uG/kyRZes
A4g9uyjSG28lOQgs8Y7E2cgAEk5/eKKxebqdonuq8zS1ps1ozvItEcW66/UQX6u1
Kyylx3YK3XCKIShvd2xCMqp1RTz8cF7nQbJuSz0yRB4mb4sTYbORKe4j9iZwNAZY
3IXZn6WWOV0zmGwANjnu03UXfhbQAY9m9Rfg8I9sPJFU7IZZflI7wCf/SmEhnc3O
eA1YixfyiNuNYrlUBU9G+9lUTM4wpTZCrmT18TkyAxaLrFZXCWxqgGpQkthg86pz
NtRewAxc4s+a/cOSVyRgOyl8DMPiY78my63V10OmYqW+Z/bY3dH35SmLkRvQiihl
LCMtVNmbmwswLanTxQD7F3tAklTcSYCG4uDFxby/IvqaWLck6DVOYEfmVptxkS77
fe1LZSRKSMMO+LXB6Z0Kj6iX32O8F9rrQBW1nnc3AQwpTzB47L7czoyA7LjnGUQS
4T3L4cyoSa8EA4DM/5tVcjp+NNIk7vSm2FiRJKx4dTWphpUIFPgfuWqVY9FKIFwX
ix/CkY4d2Lkmm/VCgxJadZTCSWnWY0vfOq4lDkOdUUjubCH99THRFPee5TT9mUu+
I0cUiNrxgSOpjVxkaYDdxIj0lZjr7A9UFPDRQ/mACOKznKK0RmMkhNA13vycC/vC
XySqpYjJ7WCM1rYVg7Z+AOJe/AsGNDauSgerV5lumJcZDhhMZMSyAEk4LErYIgzZ
AqwGheFi1FA2Lb0uUbgRILU0x58ESttcQa4065WXeL3fFS3aLnwWkqTmJtYZlUmf
bQ6CdBmtrTeQFxWgcMs+7riN2+PaRMO7c30ppyShOzf68arVyL7UwQQdnphwYehA
x8ejDQSaOHZv4F1VLPGqqlTPUrbU3H6X162frTeB7FWYEBVCS9pm7XME1eObWXx6
iHVUAL8Tzp5H0mI7j8Wyqnr14uj8+CDcZvQfTv506jTR+WNZEZDz7ydUHc9WehFj
XK7h65bwAqjHprzzsD0DuNeF+gcvAlPfvz2iEh6G1U+MnwRmkJVmjIwrCDQ2sSFw
9x2pZlgM+GDEqq381Yhc1RFGx+EbYVKo/haUMXyw0MEFW6S9J/sT/qCTJI9ovX6Y
ibsPBtSJm4zwhfiz0ygp3T4EtEOQ1O+AfNq76tIWZ6vjoHD0/JYUBb9V4CPA2CAS
YvVCnUbbch4FBnTmcrzbHtLxnDlAS2HVB4UepiYxxZDWbiZle4Z13cYiXu9WEsfJ
vzTfs3irdpPQ17FYeOsPX86MN1MubQo0qxWkntUJ/xlHOAlzaXfYtgLGYePLxptl
XAhLd5VRj2HJgZSom5o3WM+WKmEqq8u1RzR6iV23fnHu+IXU1Y8RY1WRDkOvM1ed
faCO2Ye1qJE2ZMpRKKWOfCPsYuxBaZVpy2GNBYO6NAJM+cMB/eVh4ZqYPuNJ5d4w
Q2WESs0QsK+8NX8zEhGt+I+SvCtozfH5fYG5MDo7ApdiHp5IXvDWLg2yyme95Kgi
Iflt6ecx60zRCX0gJ4MTiPTP+V/PwzB/QcJLmoF4vaLSA6FBbZ+hS96Ol5yFKfn9
iYZoB67y8dshukbGEmDYZJM3YVpgxP6+KzrMvEJDj8s7sqMuqLifB3HsA2QzoNMW
Z94jtJzhyKfk2xroGJUdEni8h2r+rssOVhF+0isX8UFd/NN6h7J0H1p6sE0qFuLP
8cxE/bt1IsVwXn0P3QStFbT1BzbBT9FvwlB9/263CFXPs0WwrkMWWW2dq8iPlr2q
Tab5KCzyBDg9lldKO8yhPo2Pdt3nGetypp1V7bd4g3KSHO6hppA47wy4TGKjESku
Q63k6dQY4X8asDoaCgNqZJ4ml7YW02/boS9xb7pdY+r4GE0uMQyV76VIWzMz2hE5
5qRSIKuhkZWOBnTSmbvU0LcG0biAKjQ9PIxlV7ks3e7q9+xId08SYaMPX1NdC6DV
rrnSq4GxLk/lc1uUP0Udx0jU5YYL3ytaUF+Vr4ZGciyEIuBem0LgAo4SvX5H/RSk
YKZCMoZLenThk4+ZRHkseMmQgcdH8cdYuXjS0UAkE/PYnWTttHerKTnlMaa/zwW3
Uyj8u5oUi8RDNBr/jwu7zo5vqOoclwUkQPDQEOR/hRmPDKMyollQpa2VfBauzMAp
1KQLLSLyYzhzi7Ue0uyW/JcrrFsem29WlykfmP8n2csTzbiZEMTAbuaD0owUeJOl
5Rw4Pc+XK1vVBSJwcD1JbEKeKgz7hrPHtaOPCo1wm+70lyFykEZ28ZmGIrCyfGVq
HaciA1qle9bTSma5Kgi+xSdXoJiEVht/pGXQj0bNjLC2UlmYsOBbl0ZQjW6VmMUX
xL9YuygzGZoyYOnqqDRC0sxen/Rl0USw0cXtSpQFxFMqV++woKs5uC/nJzTUkQjF
Masjayx/MVA9Zx1BJM+cLo6QVbjW1NNqcgBVKtyEGlRbMBQTq0Fq22ohSg0Pp/ah
ol4jDmoVciJ+qru1e/GglD+wfNK1nnlsXwe42Nj+6HQ5HnodeLlfrTjFaIbqEOrn
RPHivCh/dBqglwstU+mHKVEoLyjK7qUozXrQieNHZSUJgAF/PMbb+XfUggL7F0yW
x8nJrTamwFc06vviEQuxju8NL307uk1KijeiYGDjahJdy3QNkkNK9tniWk5531x7
ZhRVV4J3j4DANX9SdWOgj1mBCalkwP7natdQEz9teMVuhugKlSHty5CPrJ2M+J1+
9Rkguax+JyseHUqTuFQL+r4VgEyQEqeedPf/h/cYRJua6AZT2tTS+jk3a1MZBQS5
0HHaKvNogqD8tTIe0izFc65WyrcbeD/8olNKYGFbJBCFm1yb8wqfyhXOYPp+3zRo
iXwneKimZWANPwGkchxeKm5a5dkTBDJpZ33Ba/H4TvYFYCAjhrC86GgFYYh9ZKBY
i4spq914n6+ivr7g74ELwlM7FOyP2HTd5SxDafP3Tbs6WkGi+UEgaZrs4gvVXUxZ
DHomJdW2i2CD7GUni9X7hzRj/edx9q7AjMaXZ2IPUyPv9Z8bqhkJDItZWcJrt+1H
6l1L4fj3AMtIXClOI2t9Nx4yYxpRfE3WSQlnMHOmVjT9iAovj9mqYctSvME63Sm4
jcGAW3ZlDwX3o4VlnmGn20edM1u1fWWn4fp4loBW5jgPRJXnZakLviccPhCUp7gj
Edua30NSz1CGkgxTCXGcySgUAgH4Bqal7yUZtSO+ijRPy2AbumdCLaVTAU/DRsyF
CRfQ0SwfNhQikBwsF+kp9Y+k8hR0i/p1gVaYSkkL+RLPO8JnkYn7XbENHiUMleV0
kAI96otI8xRoy6J4pt1BCoBS/wIBW18U/2j+nHck2DbXHGXgbAkkLyVGSRZcAuJV
R7msz4ndGaREL9IKhK61tpbDqFFM2e95TClyP0L83SmwCb0+iCK/VA7k0IxdrlqA
t5lxjhUAP5qMWZkqEKjgpmIR+g4VJq6m4IS+TQCotWo+L2LHYfEzbifbI2t8y6Rd
qLWLKVbPk9vQ6lAu6NcixqguXBQi40oN9Hexg8IC1KnqaR4DrWMHrxYT28DAs5OV
uPUF3M6ohQrPpkcxDI55eDZHqbmSsY/fKH/HZISYdTUERlH+oiq1vu23MoU9xec3
svUMEc//CmhQBY+x26TvS0ZIICM2BFaDszoyMdcmRImTdYNsuQPz6BmWimg0/YS7
FDUSDAUguk2sK9qC7R+XEndatpgJYPtIe1Bj8xDXWG7aVsLlVMnXrXpAP3rd9LHd
eZn4mLMLNYo3QzfliEOgCCvkAzUwQUI1RQ9t9nRBK2+l4VT+hIH88wonGSaXThzC
e4QmZSxWlxKm8hOJUe+mTLlyZwdTMxvaqdCa5KBqywtgqhVoUHUGynZuh/k/c6p+
uCvD5y0TTXYTENmIm4CJj3MnZ1gi4E1aVCas+APRKB649A0C/luRLablLLN3PZNx
eWTDrjK/MMe2362Md9uzM8dS5Zh/BzunoWT44b9lGfdDZUTxC9ZY1Irebb7+vGhH
+3l9VHfjnvXoB9c1KqC8EgUUfUuz0FfYJggehuWrEVYhH626LxOw0sA0tB24Mlah
FggrLWFXH/Fw0EtdwuGTZZNxrP5UIPxE1Jume/ths/9d49gStlI/zzuBsgDlPnSM
yP8sJqjxFmNRvnPbYAIGNpZhx9eZfxeeTlKCEm9RcDW/tIwz6u4ims80b57e1LXP
eLtinycosduUBlbxZkGscTqnGJLZXENaDrZ+iJH1LTJrx3Y+eYnzpTJupx+8QsPK
s4/nu0x1AqBjMMdkJh4cOUzOOWbE41dM2iZQPaqwNZlmPmLU585t3P76cUhirfJH
yOx7Z4EElxBYByAurc5QVks1Car8EOJEWZycY2dbwBNwXSOjVI8Ax8sRlivNWYx7
AehG7g3c23fl5FUYXSGmptOw6Z2Ks0BdT+jlKcNczM8OeCT54n1INL47k/4TaRZt
dQPy5QMG8WXGOEPpI8WhvwkJzKe9E2Jc6AXWHvku9y9iJuAGpBBMFBJm72uB+e3+
1HEQOZtwBhCFg3/nmt+kzs1vQj3ucSamH+LR1+b01IKn9iM3kqKjLPJ7/MRGKVe3
iR1R2BncLmZVnUJOQYh+4Axbg+EN2R3RXV+C2WHzhtsr+p+8wca3pA55cjfBIu1P
ss6TYAsVOSqKVuVO6xbN6QvhhQ0y0zUaTbuGCtLZZ3NqQVZAALi+NV8o1DYAFUdm
hsd4Iut2+j8H7sKC2ZunJd2qO+CF6X7O6SO+jxWFyFfrsx6uXbJvRpwJNRRQ+jwD
04vRNKPW3IiKd4WI+AZ5mjgvm4Exyls7zB7BFsIO/rY1TSE/fT9CyHTAo/7AJC6A
LZmEpSaanAtGUcU4IzVwlZIkQRcdkh03xtT4u72Y0tlXKySeYXGV0r33uRcibjYE
rN3h+Sp2UHrFoyRhVICeVd64YQySQqNJSK+4+fWRwVXi6Kj0sKymS7JETkWZqzsK
VpKueWLrlBvA9opE14YVTxT9fNE2lMry9HY/Z0ABBbLxc4vgt4t3siapaBluO1M4
d/UrsvDW7/YqEIysyR5U8vkn7hdMfNRRthsk3Daa8+VlQEBOYIXHyyefqbdyo8R1
UAFlYN988E62dd3R0jv5KesWUf/MJOl1Ph72M3ppouw1XnqwIP5giQyg1DETgOzo
m72pSNtbU38VMDhqgiSPqRjIZtDd1EX2664246Y5eQ4iAG911ZqXYaHhfYGp6v3R
/4MC19HnFH7HsLHjAzjXnvbC5fpFg9dr5Yg0K/9gr8Y60QbeVCefN90eGzxQ7kTm
5uIEC8gvs5ZNJ/LZfdBDtirH2Ck09bzrhN3jqqYc/qdXM/SbLXUNUWFYt4wNAz5j
FO+ny48l1mISt4+jvtMC34wMZzoM41WHMsuSbZwLw8hjCXauiaX7JxLO07oL+szL
q37qBfwcvZOzRNz0klsCAg0ett0Nz1/LWL8UWMvqdb0jJF+grVrPCB0WnigRWKLk
JD/NQS6Nqn+ytf7k5cNMgzESn1h8SQIrXw0XNmc+1Pr6hATVAfCwt+Ofqspc4Fl0
4WTxjkokcUi1WRsrmdzVwuCiB3aVWTgE3d2SFIidNlEcELLecAq3TIGHeEcD6Eh9
qxfxy27xhRk6bbdwnvOybU+A6UgWlp1d8GUNe1MV3XcBYRfJfocXHIEugBMpVGQb
/rt808qUQV9R6IwVixYEHhukkEZ+2tr5VYExwurXks1N96FVA9LHBtT3knKQ3mNN
ciRQdIPGCkyMkVpN82fAHGUSiCYcTUXacP0S8BWPYF9dnM2NMdC0VGfjI+uvf1nH
DsnNnjEnFjf2KLynzKQTetfLsGCmh1gbehA+lVTOGcUODH5unGRf/H6PIsmrPKu3
8e6hddmHyi9QMt4ZnWmhIkMLI/lphEKUvb90XyWp+EnHeFDKYKhbibo+8/NZe0ez
o6wUizCNjLGL+XBIPbx0/glqExeibQnrHHobZCM1k0oRo9ecQmyv4xvMfXry2EdZ
GgvBuaJbbfvMdLcMN11yUtJuTl4fJ5Mvr6vSkWvxC+B6mAewxKol0Kx34IC+ojOh
SZP4Lb1LiJF8rqNlR8ppe9P06C2K7JEx0J9C+hMOdsX6cQiXzghhb/FdOQZM5j4m
lYFnCvO/giVyHawWfzFwGcSAgsfGSDgY59uz6it6x2rN0NgvMKAGcphe88kPfxlu
K44opZqMvJxcWSg+jUAvwdxjxr2+4Q9JTfLLWRQvohOqjpdO18/tFFRtWchs5Gmx
A2y1lg4hrlSJ6EoukmBiwsgTBpWwk1dEabrsiavGeHHN6B/ER0ZK9Gq0ZobM3q3Z
UY+l7nXI7jaVQFMxI6Hji5w0YCe7jlpqSLWmCCJ6I8b2lBmEYv8qlrR+BFx3rrLQ
gKo/zRZGyXhDIxPycDQhW9MHZCCB2BwCUU2kwLeVwmhd4ZSoPH/MT9HSRr4sFrQJ
BI0ZSfcZfhK+6gHF1Jke9f4aL3AXvfzgSO+4DUPjDRZp/yxIqor8ZG1m6Mnhdas/
gwuSmsNymuxEc3PDuz7JX+3gs0cv4AQ2IMtZ99h6EhTQk2RzplMo4/2VbUe+6tx0
mOvrTt0JLs7WSzfOkxUJGFwHis9xFESdYlLn2j3ST2EfziJ5s5pVzybylRWRZJSG
sxFB/NB8UJ/4BkYbHcQCK72OR1efXqRLfBlelsKPj3I/4PHMUgZsokklXcBmJcvP
mRTIi9/ZR/SmPAbgQ6Gzh+3XmDXOb0rdpsXoNGOhzwAu87XtHSjPhOq62vYUJpKR
L9oogyAYw91F34AaMKyIo2YoylwhUwRSHcGVimOPxGE1upWQqZN0L2ElcIe543Uy
pEKKhDm0BTCniTxNKXRleeWHOTnWviMOb3q2xeozeJNDW/5k9oygHYVLjozshbyp
2mTSUXax0/LK3vg6p4u2FTjYH5C2Fn1CPK/p7U0lf4FQTzHkgiCSm8tbwDSoBAGj
SjSqfvkBEKDCF0HbBMVqBXTOVuthiphiNTejFRLJiCatcIZuloBR60H2BTnp8aVn
It5hREQf0VThDE3lUIWNJwTEzWu2sZtnMIffxmW0AuLPaTC9xhnv+NXJKJ/9ozgG
ClE1+Mm9+lakxPT/jsbF/KFBpmQGU9Xa/NAZN1QdbUAYWbiQzf4zPT6aXym8dlj7
+82O2EwevJPHBbD7OxL/RvMGGPD+hD7SjNWNQ1yYmk6rDxMI4lZRUkDUarFnI2Gu
ghUO/d9A7DhKWFw7McKEKNDwyez65mxIKGn7TDmbh6yli5kr87T+Dn8STlLmAwU2
sEaVBg4yBqY1MVlYLYyxcNz7JKcdSHQVoRJ3mYN25lx5W26YAxJ+wUWBkwKS3HrS
9ol7jR5TYWzdJr1kIDk/pCWRbO74Sb67Jw9icO+uNW/y2OSAX0L3j/ef6h4IGGfF
T1Id2ySZvPWxseDc5Shm1OGVlKky6dlwdNcrF4EtFW681jXNbNDoOliMpgOHdor8
bFFjSwZ43dZYxHbhq2sYtunoekj1iK79qXopNPbZibJYc38fLw0l2mb0dao3mhs8
h1LLU5BKBAxwSvs3WqDzwcNT7qplxt7FnpyWOAkWFjRMA4NESa6bieNyBx8tbZ3a
AQ9oH9A0V8pe2pBF+jTGDhjPcIv/YoTsgh+pZ98ljrFTUn/26U2gd8GD5v8zyWVy
RQ6HIzGHmmHz/x60CUNWl5J5xXwVSAbRkSi7Nk82tffwYE1RgCrRvym69r6UZXzF
nimHOyysEwXp/jXVFFTntTSeL5ZFvIoMKgTYT6xZOPUQhxgi7QuuucLLrexjGgKQ
n1eoE26iLMHqfYDLM/Ok4Dq2tVOfSJu3dmwbuGB1nKbt0NquEwB0lGKkT7b2QR3S
gg0mFRuAkNNA9DOZPWnnm5vH8WnWrj5bQQ5iahtJ1qS4e7W6+2vYGmpZZQbTZG7N
1FnN00ziObYtBjEsCIeLxHLcdoT5UuCDYFV8TQnwKnGD1X1HQVkCZHC9x0KasUzA
NqYGRplKzZBoHlA44LHAuNUolH4odYnFwkXkugkc2xF73hdp7c7kEbx5gihv721m
xR+y+EncQ0o+ZHHHEykHXsmp6+Ey7X4l/hySOJM2dchUFW1DyPhqjU7LdVUpt8dR
wAp8GkzOo0xr4yC3XjE+3hIpYPtVvHsNDO+tTl1KsMRYrON172rjxeM1n58VApYV
4CCLhBQafuFs4ZAUXXk4PaxOn1FX2/+qA+801yBh4hlmtBCI95iH6JPgJn3Cy+5u
6tw1JovE7e/2GuLt1uZA5v78EmKNLZ8auMw3mqx0QkBJE2f5OJm8Il1icFcnfoX2
1cUzwWrBe8S3tnF0PkvtTE58+CUq0b7rjpspV75gx7kFxZMCp8Bldf02t58qGxfV
5cMdxxPxwuKhWV/57p6wRpXblv0vXLQBzPRkTUuIMcgcqim1trwLFh+crqtsBNt+
b+O34VSh4xgB8DPlkUgU+6UMD+FBpzTj9jMOcAOhD4/g3Sl3TrLWybapYDecDm8l
kRysoXER+VdCeaI/48x5wAvAz6avzzTitiY3qddHNgqZqOleiJz63aOn78k10CmC
kcPIvZsQmFMewTg3mqCTJsEw5UMhEAj10yC7niTmUDk1Zs5PU8WlCaToxO+IULQZ
rIjRbajoc4CgqXlC4ZI4bHnIUxkGVOOdGCMfzAviR+G8r6uAkBI6O1lxQthvGtwO
wWopZMrEkjFaMPQEcNNJOYIAEnRth4cfJHocJn507le6YqzV6YiapCW4d/yDpNSc
3lWJwaxjweLmGJNNhqqog4RSaNQM8fU9jCZqdgVraIxd1w0uy/EmganlePpWrlEX
31TJdtycx4POdVHRM4FRl2Je4oBvjQG2KeHnfW3xUFPrHht+fa9mYczvqVBOViRw
X7rIaUzKX8gWJZ8UVYHfv5eJ5CsAqDMScY0tWL6XXH8r77oRmzw9dJBQggsTiu/1
9+px71rMCHc4UCIQiq/+cq+Kut8SQx8JNEDuKDjvj2U8/iZq2vUt8DFlDxfbd2tM
EzuomRAP6rt74cFARsX/H/T8aUWcqFspD4WmQV2zazVvaU6yioY0SynA3FqynZbv
1G3hbdnW2Zpt7iMOEb3W3ujI4frfqSrZSF880q2lS3Bp0lLi1Qn5brZvrzQhaOtv
IHVkRL2s6bEDnKYcCuPE6UxW1+5Zc/DQp5bmEeisjm39aaJqJpaOQ/5LVJsmo4dc
7XR/JZRWu9nipvAcE5/bqL8EKczchO0RHwagNP5DQkMocStKVE1fth0gvq1bY6p6
40WvmEMwSei87LskmdoDy/PYrD+T2r6Ixo7hU5WbrY1jh9Rcie8BhN4j25IEQXkw
Yb3pTUNnCG4jVxXzFaTPAD+OuJ/Xrm4NvC/YWOG1OBTLv2bo5TNVmf7eBjGZ4dq2
SuqWf6q7i4j/xKr0dZD8aRvlFPGs3VL0yZG6mWsqOcdpVRcA+/MCRY2XQp9AKDKL
3Wz2es09NGmi0Mx3OJXhil3jJc4Bl1RMOeFWxjldCXdpWxJbrTqi3ZuUARoXYioU
WrRyUwcKo40usRnKs8P22NxTNqTTScQIWh80zqBeiPFbNTGaI0VWqVTL65F3uUKs
y11HnoCTMkZ3D/yFkFtKKCAogPbU0xj3fwWd7artR3Yk0hzBJCcK4iWUIaplc9A1
Ji/qARn71bDLL7zKriqcnQEQRCgIS4DwWDPKmRwEDnjJ5dyh/jPGglyqpBeh/gWh
H+gNw3GKPnlI3iCxevfVNhP+Sv4xedjyM56tS0aSs9goudXIPFvugXgLo+F355yk
OKZsxlHdwijNMm5EVwtrr3/pkOpwU2Uu0xfDsqPKPLUYWNCmYjECcN1ojGb5YNEk
2wCLkuycZjAA6tByspuNyuLufYV6KFfqXpWW/le1ENzufYJlW1dpCrN3Y0SUv8BW
BjqA1Kc7IpMlqZNcWQh/9tKhMfXhL+3pWhLKHRvuJbm8R2uv0ZpTk7ZEapUZ0TmN
iHlLYet65ySNx4ai0O5dxbpcetX+OmXmZqKabiSks29Cc4Pmjq+nW/md5c8e/SD+
U4KqvR9p/8tcIfp4NeEmZYkTLaJd+i6WJg82za3y18Dxb7lvxtIgNLWwE0vzKcBO
uM5cYtBJPK5RCJ6J89vTyMzifGPjVlpWbGD6o4p9QZdoAlTLj5u0lSfFOOd/vB8I
J6LHWLtLpo/VXQZ5enrYfqNvzeyj1Mf5+7USM+dNCAm30zLFginyU5ZCeO3hK692
RwEu46lVHMZKjLThvBwQicQpMpT7glpR5XHKAyb47VcuY/INg8YlvBLcjii7emLf
/zCjFtOifIaAFpcgA9ovXi0vnKj328vSyAsD5lN7SGUHs2d+7A52Zsa4aWxNmAqB
8iFakOCEzzfkUsBpzSRvTQ/Ju/RDTCaU2vRIta1gaLzLcz1oUHLN4JU5DdxxlfMq
hD/jQU7CFhTaxPBBbqm9moI+wxLLzQTvs3urczZ3WuTRtk5geoI53ob2o1VNsAh/
ZRNrGGuIcVDy3kmTbU9EEFYwY3WDGFH4vkyAaCvfVq+ZxekeVPQpDwMr2DOoqMtz
8qQiTTI9rlMZ9W9f4jl/FYdT19qKAha5nVJiYRfN8c7GreazzuMB7eQlo1gheFYM
K8GcIPxexysRe0k0agjmeB8jhv4pANSTuKbwd/0XaROngaocY9pcth8Ab/L+Ppla
UIy7ToMayAe10W3TgBDXDY/w6HPysu23jisO8rO1xJL5/3DqATLeQXvAgWHgs5OO
euEF2VASgodF6XZBPmycftAtvMJ3IIsx7YKe0AkdMU/gfgDhDNDPiTMgz1zxioF/
iEuwi/iQI9baDUhNA1mCMk8M67cqBwqzhfANbEXHN6oeiC+5lDCKBAjXvjXbq6+8
LyMOS0lPW1/rLTY/OumlMHao+20bzcF4A0aDVSbB5RTxgLs9mBr3RYbJHv5+/oBN
3fwyWrB0Qzkdy7V/C1/9RIkM0dJlPHVvzU4+Ksfa1tpi0s52ru4rJUUafkIoJVkD
wZLgbpstkVUx8W3yqvH9xXfPG3Z88uQZIcVE5+GcyJ2SdbUNl1kDwyg0Ea2McDYZ
PzadzXV4h2UuL6MUenzHz6dS9IZXi8aNP/2Iw5PDV5RH7pW44j240DXlMe+A0NTQ
w1yoCljzZ6y1G/np62YbSZ1VkOKoQrR842GwWAWmgCDO8hIpxs3RByivn8Scijl9
L2T3FSIhckURdrkM8ieWrDc5KFd6fRQ+0aBEofKhPObs9YOvt12Au1zrfkkMF0nM
DirjdKFtmymYjL62NAsc3ESGJQdWjuwFFHa0UClyKSveCnwnoGuZ0QS3zWjXeEsS
+pFIp5lgCCzW1qPO2+3oRetnRupBzLASLRD+OSPMYFjMAur2044G6Cox7zVk7x0t
tNM19R/S+0BD0ihWwXWDzFLVYQxM/7T7WhjbSPvgMtWuAk0Y7yecJB9/WLM0ct1F
lwmv51367K0gLFUqVz8nsKZkgtVvos5rYMwxX/j/NQrhE/2dvrPmrm2cXrZSnw02
kyemCJ6U6S79aWVHDkNu49zOIMSUe4IKrstT+xRca2g2Ox0bWD0GKWbqOkMGFrtK
gggIeRzxWJLajL1HXewhpg5yUn9oVXOJTwksZBMmxKmnJzKC0s9m8rZt+D6BQhiP
nPiAhVwv2NelnlzvkN5MEdhWSAdQwfPJJMJwSGKmt8HbT5zz9iEkjEErEIvzyQI1
N/Heq7VWj39AMELxec/SBO3rRvvg5pOU7eIvCZEiFIwA2PJv5AsOLxydF8J8bbxI
molOxzONcfwLwCIM3ixy3hIxzdVvVljoAzvlzP75UgVi6y5SDLdBtWO11xBjYAqo
R96EdKsL0tYiX45vVJWjbZSVhoh6HDj4PhF2r8GcBhkG3yv61AHzhK/ZFaTVyp3x
ZbMC34wc6NlbW8cwb//uRtQr+zvTeLVu7Q8k0/Suees8dSYIBLonR5GKN07GQ18Z
swj4KUfflR/yZxzXrdKdYFjM8MyM6uS63VLcghjuqC1QQmwp3qy3yhKm/gjMph8Z
bH1uEw5ceCBTVMyj6QLqBLBFkqnneQw/sb7xgValepqL8DeXKoeN5CxlRp0EEyCV
GqXoS9zVh+DZ7w5YupqbacHQL7Xcx8gAdJNlIwk4WvGho7swKjcEA06/oaPwCZaW
kX/k830cFh8i4PyamJ3TKx7nRorNcdrI7k11bEHy6Xuz05bdV0WSEHmxYYVr/JP9
EsSyKKeVfsRcGHuiKBbA3/bWizk1bRnikHH4ibzsNjNs86xenBrIYfgHWDuZ4HCu
mcaBLnNjjbmDq5PFedjMcJAV3U/2j1lbNQ3zBDEO6o+RV+LsyiOro7E9FfBsephW
wbJPw48QmUpiVTIaKcFSuvQLca4Gm2D4tdiEbRehyShWXtVCzjT1OJAhzgY6Q3Li
KAZ90TD475cYy80EkRtrcs57NHfVXd0oc9Yt9fcqD2qp1PDkZnsYYGDWNSSgHDWP
DYu3Euw/MdvkJxL0REKb4PG5Gdw4iiEM3pWIO0ST2btQyPQmkh9ZI5ZEYLwnSw+h
qTumItEHLMjQnjk9ktKWutoDPQs8/lUC0SEhPEwzq+5fuFzP5SVvUXeEAfVeznpk
oM3cgjizyksf82YvdjwcE44HHSTR64zIXelRpYEhAiXarWhnOcpm1QbxeExUZ2Bb
Af5e8L1bxA7hHtdF2xh9UtnnLYG5WuWnA6iCNzUVuE7pndGf7iyHwYGt/q7zbqIP
APYBG1/3enuJkPfkLqwzXGklHKFC9pt0GIcHHrB0iwOP+si54LoK6ShtdVhOLyBz
9AppCGzIqJyqite2j6uvr/ZNp3gsTVzQlY0A88fIgd/ivMZg48N+pWnTJwBa/dIj
kcFFXGHcW6PNjJgbERbR+BVa84p6T10I/Wr7AldTQHAlzoG3RUPVCwYSXS8cO6ZN
Miisam8am0RDvlzZwnivQhu1HF78YlxY6PVEuRS9Dn58koGQqn5Ad6dUGUXl4BHO
SoF5RSCIMD+zp/n2I4KJkguE19Hqxl5qXOXMh6/6FRHTT2ykmmqAUrBa6oyKiDPm
+9e09WWU+6Rq4dNkt5ELb4LQLroNaPU8wYbTOXHCNFiRVTtM6WEJEzNELNzfMVjj
T2lwlg8Je30tk7d9BTlRnLjYF8NJ2JEGksz8xA8gfH97n8HBXWrKMWo5tQqKcKke
ItztgFn68S1sCSlywtjhfBxduvL2qL5ijqUSYa+xzViUPcgIuwxw3Qww40jZDDyc
vkk/ZQKCOazz930EXyHJpq8w/iuRiEjKbzEa0+ML4nU5WfDtNoAuZ0rBwuEFPMqp
c3EMjcvo30YHHWm33b6uaIPCIJGNOsS/yu/kf75UlKg2bvRLTn+zXdPiizMJLyk8
bgNlxLFVnR41kCfgd0I+byhmPfezZqFY2WJAj6nGPU28ir9Japqh3ACpqc0GdfBE
B/iN4H7Nn2zIlBJdNHINCIZqcFsMfat/fV37F3cX2F48D4yYNGIve9Hul4cX088f
piKKKrk9ny7/6YCDQJuTsDNM4dY0/1s+KlYp/YYDZofEurYa5cVkJPnR8okPUAES
HbMPqtBILPjgNqYOzOszcGsNDEeLA60VmNGNa4j9GfDVvEOjsFA5mPdAN4YbMsjf
Pj6+hVVFBxPDgGWgTRZsMz7gdmTMNjtm9/sEbFH2sxA0jUp+wiLElst1QzTOpb+r
GUmvDog0QyQrmqFbQyQar6exLgEtA4gnxRjBnTVt6ydjuK9pI0KUHL2gGwGdGYp7
cAXVjcB/LoQWSbG5b3t+8vF6j5LxASSa1Ta+p1SGjDXqaDuZt3nN2O4pDA/jN/+t
sIdJE6qY1KuPPksVoR417H37tgKj5rTOBdJXyX+Qe7lyL4yWJNYBahlzQ/VDUmHw
ibP9BJMZzXpI5t5hdbYMy5BjFIIQteVg0l+NNQ6jHqFAxkpbrUL0kIQgG/kwjZOw
VIhdW7qz+SqJCueD/5VdcCQcmbETss5q4JWH7B9SISRcx1VH7z55YVfhgiMIYGtz
5JlP7Dbd1P19yThLZyLbU279u55xiPA4yTwewoj4l0sqZ/aPvKHP3ls+IdBMdONf
zWttmqnTly6XeXWtIyIyDljKDEW8GL5y0wUWSGNgdbshIrxx1ZjnKwVI82Znh4td
TeZxN1i9/wtYWv/7/BxnrrTrZuGvZudWwenSjo8y/+uZ7P9kvFmb7BXgQrkXbFV6
+2z66IC09mX4Xn1tFM9/Mrf+itNUyHfNFXIbdEomdTV4HYb2dJt86pVVjVQaaBTi
rQFYSTH2ImZJE0HiVrsqQzZKVQIlYbpkkDeKpSczgAjIZtHuoSf6TftvX68u4RZr
YT3vkv1wXPZpTjU2/T6VS7fpmBm0c0jWTD52if7AkVbX3cfoOuweCdDFAkcd04XJ
SOfOMK10sOCYZu3kj7cGTPrMRTYbOYN4FSJwHU1FHq6rHSUxORk2sP/U1eakDvLK
56wWKD/7vPQJCTXokCUKBNMt8OHwSguYtggjfzl6QDeZsllzV/FVdzJGrstaRnzq
Rv/gOeIdDoSoRr/iFy26QC/0D2haujlDPFH3rY/LNuVEDctw6cBELUFha1HFtkRn
cwfQJeFvLeSSulnbjofMEvyuDNxT6pQF7zdJDkA+k2l5IHS22qJa44Hzb/iVyHSd
czCF9wgFJREhBSyPGIh9YeZdnJGb/seRNSsdDbKGo/MnoQl9VK85kMhqz+3Zngfr
3zVBGGLKId/Qy4vpXlWVvhc6GWEHLzZ7ENggZOMFR4iM79STzCuDAtpRfAknq6FS
kCRKBBbwW1xtvWEqIAl+2JFQCtDh5Ej5sl2iTJ66T7c+RMRvHgwetlcNGXWHGIHs
stmIYO/FM0U0jVLBaPjrIxDixqzDlnh+yn4WW19A7S3uKK18dRb34ksTodKRiM+U
NzTCWYZmh8HfPU8BBHNHyZRW6FQ9eltMDwk65wBnMFA//njs2kFdVlcikQCJaz1o
eve+eBZJ7IVMBUKR4TyDP9+SkE6cEgxeMfbAEDx0Yk3dYpVrKWUDpIt/zGk7N95s
gy7+m6NKXsZLGIvvmCic+CAGMkP3ehJZWuTbnylQvtBTBaDPsCr5hFvZHtHPuzY0
fLrDsRXAINUni29iK5eGdxIaz99UBo7zlsrv+SRSPFzZ4HefW6F1O1jRzE1hYbhE
/sj+cGTMwwDRzQtJJPIfUmFfBtoQJkq+UBfe0h57U6QePikMFKkbt1mCoxZFvcMy
nkBYX/BfA2GTzfFuqxhw32TbbAU9vT5P9vroy1xwUzudX//U85X6iD4n1pbvpBlU
b8v1yC4w5yY9dfOI+GsrwZvCT4KYfUT5rkepkGa2/6LyNgh3fkz1bKyM+cJXP2hV
v4qBwlCevGp3GXYMsfTMregWRoOx8imBu4yDxWC8pZZLUagv2P+AgU7Xr8SyMOat
TqE5clTVQxG+qtJxT7ueIILQhPPp0R48R61r0Km6FUPEgziTE1AEVKuoP3fp5GrP
fTd8GtPwdaX6PjkmDp24RnUauMft5fzS851t1WZWXr/ngY0Lnao2KXjHUcUHGjLY
euuHmplDfm4te1sqFY88svz28MOpD4zGWWOv9yalsZ70BzWbqIYvhlJCxidvfNtk
VTmtE8O6rWqjB773whfAH968L/KOkk/A719WFANL0A0ZVN/ShZck5y7gkgp20x+z
qPPVtWqBivlKGfdHAr/W5FBoXIGX7cYBVynVMEDBI1sA23GMNzNzw/umYhM0Cmse
sh7Y2Hb1usExyIAElrzhLy87lwepSZqyDpD7/8q74VYXSPGtT9Nn2SM+mcghtc/D
hGfXj3yQm+oWyGpazGmOQslOo0n50apUbj9SeX/l5ft6kCURwSqEEWQoHmi42g3z
EW48DTpCtqnrTssy9lvUwTm5eUE9TkGLBHvq3Lzfta2U/8R5OixL1J5frDtvRg+m
gJBwL0vLCopOVUWQovAGjxfkobV+I9EJM8rihasNmOLtiwIBKNlNtTf/chu0be3K
5dnStvIvCiNtvQk9fdCN626dSLK2MXF+wnsxKP/+h4F3yGFOHjLIMunHbZGat3iF
zdrlQARy8ZAinDbGhC64HDJkuCsEdPYaFSjJ7OLlK8UZhBjlUBOJukSp1CFSnwXY
TaSz8z1uBwBN43f4y2OlYuLCGmk3LeMaxhUFVYvs/qU8Jk80gR/ZbJ6d/PDG5smE
wyLCd6HzaVvfgimSuiKx5vLpEFtTd6lZcw21sgfHmtgFjs1KAd9lAJn87kWjtySn
fskeVuiuRPFgUzGr8S5oQUHRdTq2IuMVb820HcY5ea/Z9iK7lh0AtDhqLA3uxzxm
/fB22EnVD4LlCjPS5fLUbQzxxsxJN1UjqSnqlgly0ByKVPCwytDXfk8frBnPSidK
ge40vpgOez/CcYN4IHoRRK8npYLKWGqxEHPE3B/DOQGHHDaodbVM3FKwoEHUCT8F
mxbVpNk2FUtIiiiIC3pKDBj6tk0dkbmWyix94NICKxoceVNi+z6TucpRuDP7ec5Y
WvpwFFhLeK+o1omDRHnV6xTOpN12cO4RYQhI4QwV/qBvPvOKJAxKjfUzIzUlU0sn
AaGe3N7Vi14oC4Avrkb0s3SnClg8ZMFaM99MvGjCxuyy9ERQQh1Kg0u++ICQkjl+
wlHg8h+o13Suff/mwxusrP9hPah+RS9FuPTyRGNdBkQ3Ttztsmdz127qcbQIfDrZ
aKiNpCry9zVjd4Oig4F+S4jPQt0tE5MBvwCMy1sfFEeQEW4W91vaYv7nLwjJTPfs
yhSMts/qsohF4WL9N1GIKn7LqqlufxEx1oj7eJHkK8ozAzX1It94FqtwDOLmHLYu
rnfySo8+nF6CbAMb6Ibjxq94OCxBccfCW2QBD1k/h7SJElBEsdEpZjn7qu2/TJnC
0Wcndf1LFEtLRr8b5GFCGtdHTZdqEe5q81HSzDFmT4XICUQNSn/lQsyMdWX0zzF5
5WF+IcgU25tuD9YASXc7HgOy8j2WFJY4thowaOE99zmlpBOlhAinKe2HDX36ePtz
jpaDXYwBBJU4OFmWvgsp+lKUHkvGlKoQd3TVhnbltU1UoCb4GHwUYARm/hAjdt6l
a9ovm+vE6y9hHfECQUgPV+JL2GeVlz41jhSiI5wrlBXTf93mrnHm6D4QEMWno/Ib
bF4p3KhzIeETCebR1VnLkHsSFmy6s/i6PF5S+5WWB+eAn1G0fGyZf/cFdUZH1GFC
ldGIUBOR9UCM+I8+XZDFGUyiwHneULghoR/KV6WL+zWrbOIxJotBKgxe0rNMW7oZ
neoJ7D3URAHqYuhaqsoveHQwx8gcnAzIZbMvnbDmnFekUjtRNWTOyrELR35Y2omE
SiFjk37DoFCvxppewenubXKJqZEiA2yU4BB2J9m31JFEUQnrKOZZ3pkiTBbsV7fP
Xv3aShN0pY51Zh5ur6iY6IkScHpPYB/pFCIZZAJ4kdSLuWP+k57ugvcRbkDneEEG
40JKzSHaufg0uj/tYXYJHnUWpStNMtNQwo7oDvF0KeE6y5iz0taBcyxZ1ZYDEmXY
YOAsAP/95Zdio4bK8T6GWm/SIK9gn/X87I+VdhXuNEw/VAiPk+Q5CFVwrk4W+p2W
AiFPKFdl7LfdeR4VzONW15bPt5DeIyZTxjlF2GGPVehpNSOpCCKpxPNc3XtfUmvX
bc17yTfN1SLqSgpA7Vb6WpnyW/gPx6NsRYyBN6iuIw0NVw2fgjr2OozzJ0ljUihi
zcM1x9C5qqXfawYkpPQrGchTJ+E374PF8GJhQvBmpkBoF6WvLTt2dMr7TVJsk/vn
Lt9I9X6F+HnloSykpZdfMsmmjuC5Ru6NDjqzNMUS0kZDG5kcAgrBDQupesN8hift
dGsZitqUPH3qB8RGjpfawOTXHuzl27rz/e+DRWCWKomzh+/yxqNI+H06puM+jNKT
u5xCmHyvUIv2WMAGgKfHTjBsHBKk6rMW2zvaVIhJNDHj1z/d3CWZlAx5v2TvwNd+
6SwN+frt7ygU/zHYWh6eyYDTofkMNYPquCYYrtfSnxWnyTWa10lmkbfnmig/6hbd
izFglygDMvOIgediiM828V+OAkyDDmIlVUYNianYDz39L0b77IbZ+MdRz3nEmirW
d2C8PKGIRqhs8mEDH/ZzaDHbsOEdcVgU2CzPNR5oig8yc0i638Egcu831SW1Lop0
W+qf+pwnioHGWv7UIyl0cDMcrJGy5rMrrm7e2JoPyhObrcpkbiBjMxl35tiJ/aM3
yIJpdd0gYPh7v/VzRKlYQZIzQTlfLemE9tMwUsr1dndTtyEL98Q+sUQBAZBzVzjt
NyMKAYQ/u+69b60qsWSyMlZc3gKoeFa9j/wdfrvybULRDbIpzeihDDnfdg+3C9Oe
oYJI5RiiYFSUjSPiWMqwS0qhq76e81/XvwNIHjkikPXSqwxRPA34d0WnAkJT9Qvq
lVwBGNJJl3QKdYtYHLubIWmeKFmOzqfd484VfL4eX6Ni645qtLX8MzEX/ARKSPd9
MKqHGSacSqGvuuNj0GN/i4YycVuSE7iT6GB7mJytnDcywzO+plcQ9zXuYOOBosmL
PirB+E1MorI3/5rPC5dnwolWIrKB9ZyJ069p5vLKKWb8q02ToZgd8MVHnytics8n
hQNb5F9rdAro1zbwMZx3sjcXkE42O3eKc5jmjWHDJTvKK1UapdUQQSYuc763EYry
DOIXwG/MdHb3s0wWuHpf2hxnKCQ34/8289dwlCBApGPXMpPZdW0ArG2EAXog7BQy
dWQqene4z/tiRhTW6n9zdBgLEVkPQKSek2YxI1BMUzXPFBWtoEoqUuP1pvrARaMp
T9mTdQAhbBwdUEZEwLyvURfRFlSSO0Jj372Bzwn13nzdehIS9Tp94XWedNZoQTCF
SGTMwCgyk4jGI9CgtAsaHVXSy6P3Z1ShY0JqSQRv0NSXhgxUeMxXCqmAT48jY3Kc
/7V5twzTLaRH3q6D9vw6Y8H2eEOLnB45nbTHlYKergi1FTfb7f/zhPLM3sPVmW/B
zjTLAXjatmTaGfFn+NhdDRxn2VhebrR/bBWxImt2T8BS+2pAn4yfDVPiWAC/m6ou
yEv2xJQ0htRJzjHJy/em198IqF77XfJHtVUxhNXj8u0uNR6qLLoVZBp3PxrIChm/
7FKLgmrP07414Mi7CbmrlgPmQRG95nPVZfb5IrJQzJ0CCTUbIdEsWAp9Nj4LdSbu
8g+bqvPkR8qWHxdaTsMZkqnTN1ysNzq+2ztV6lEWCetg1kUNcrDFS+IEuCfr6Eey
oGx/aM1+HXILixJtbgzF7a4CmxmNBftEe/GEjp5jgI76Yt13D68c0+Lx5RsQa30q
qI+vGw1qMuQXe4JZpFdn5d9z9Y/3XpKjIdZkgF+mlOqHTWdoxi0LqRemsr3zLQnp
JazgIvf/pQlh8W8w+SSyMoS7FEPXX5qTLZuoJppv97Qwretu05yVEAOOxgwv9VjP
45iBF//Od8m7bBo8quJcoarl3j+9YugeXsuT7mq3avo8OSjpgJkqZq4KTPNU3GXA
7ewlD4nrdFTmk1LX97X26LlkQSMBA6eNkb4i1y8CeUDj2LHIVFInrJ7M0gTKcER+
+y2yedI22h+/MGRPPSggbhZIotr/MWcvOMHel71VYnqXnmOk4GgE7aXWwPGZWUte
P/iO5AAy/NirC7gF8W7E8npixf/EfjXRTbMWBaWbrx3RdvV2e9/dwLOBUhdYR3yi
1ME0QSn2zG6MmlussNc0qdOpWeR5TZZSaRinutNKi2+Xb55LHGUGo1dBTuPtDTcC
e7u/wEZhPjglRBcHv3FOC1OPiYt0lAvI1vQ3VFz8HiuOgmmM/nJVG8l2u3n+Zsps
7BQNDyIBrO8OntXn44L2tEqqEGIM1lK5E87+gavUrQys0LBQ+Grh8mZYbtpAeCNg
9rSRECNTA81eGxclDiwcL+nHsXW5JvLjgyv5LrB73cENHRydy15/Pclolb8umIZ8
LClOe+IB4+Uu9b/akjBfpN9oQwT3DY+4mytTUCSi7OajQ4SNmzdidiGM/Ng3YvJl
tzqRiac84Tc7oUEuMvs/hH63u36N++BApv4j8PD/sVquW9b5ONQcGmy5m+6iyOb+
HFNf9BFlPxrDUw7TmVdBSP443hhbAt7DyKFXXXsQDueGmGkD81n0rhnLFciOuyyE
Kr/T8zLmkAfkAy3BXvre3fTrhECDSm4EPeWyCoS71XXbf2x2gXNwA2RDSmoFh+0D
P6GwKfum2KCE7lM6lHP/XD53bbdFvV7ZWEci3Bzm/T5EuGwS4DEv6pQ5XkAIsTQV
SsXoUuUsEW50axRs1QNeClMg8d1v174UaNYcVvD/c4VoheasPJ+mPunVSwkewWu2
S2uyuAB4WuwNr+4LQ0uQ+Ey/aHjiSMFXK2Pv+Z8ZW18lbHPx/qHp7v1ju8itCect
I1KO73OQxlBGHj3B5jTG7Si6WTvYJify+kDG0/X4zbPlvZQRwQsUCMmlcWObv89A
B20kwSB9DCr213nRQS35yHaUXGxfy3c3lr12M5WGC8Kc4S0RyLfU9k9zm0WDF5Cm
HrhQCEykH6H0y2kIbWcJMAeRSDf2bU0QDBr1g/u6fbQSFxVhBGbgsqJKfwe3H8AN
g0suiUjDpMWwjZhfUNNeBmZN0Z4XCyPaMeBQbDkqHq0t/MG8WownDjO0z8J8nB9M
qx8G808CYTvQ88EQe9eNtch3YNE/B+yy8qD2WxgR/Uuxnv5RY+UND2JKDumINI3R
p1LDB/zN/YZpmN4X1+oMMC+y2NaSWqkOeXyBEUzKAYVnBVwbPTdYe+80bQzbWyB/
FeiFqcyu7svKNYwfUf1ZsUKPrVmnDtzKNo+Tsm/ti/SWNdbbbZn9fQvuHJtrZ162
kypSF+r0SVWcNneSADfPMlM/183M0FWg7MC6560i6NwyHnG/SbExWnwPJ01k2ye5
xgArx9idvr6vnGD5oAwGcx3kQ0G1E24EajWI24AneL/wFj/OH9SCxdXvidnIQIZM
a/gyKx61KP3KCZvmSlWTAgrQu5BRnD2T/ZjD4wbrE3YDvk1+/Pf5kZs3H+OM/1an
CGj516NWeb4Yj5ZvpcF+x9vdYE8Se5PN55b1CrzWpBnobHeCS7u2DCPUrr35/Qz+
miiY9iECSOuiszMI9r3ur4BAwu5BFkqDNjUI4J77Dfh4mYfVwkKKjz/LGVM80f8+
0xXGVFzKpt0FuAz7mMm+CfzknyM6HJkkjML7Kf/XLAUR/hYHL+bgzUnoWeVrz7Xe
2u9hQtAHOPTeohBj5/esHyHoFB336Qomv8zoMakPjiWIQ5CUPt9Tou3w9HLgnzCR
3cprpT4DzR1BbpJbcMjGQeZWwAnKMw47Y3n8KAh7S25oBtX2XuUzbTL6X2hz3n/V
IoXiPKYXnPAgSEaTyyxLYiOBEZiPTa4qijk2hPZYQZIagq9g0WczQcIfxM03NIwn
oMmQIoe5mjo/8gdBKbUcxmTdXP3xDimjQ34nb59gltjFvGCBJoJB+eTr7xgIBpbR
koVQ4i9L2TA1rvJ0Y0zHFoMQqcDJ+6D3ZbsXe0VZJUpOng304aDWEeP0Nxhs9K/M
o6bOlKlT5eZw3I0YvYqlF/p1pXZSNLsQOSYSmTOb0odGdo8Lra0LgmqZcXlM7j4r
f54R4uI9pmuJQK48zwVGlQpQxeCxhpJeUct9H1dnikUxXBc/NyvjtAhlHpcppZPy
Jbir0mRfLf6s1VXi32KWRxfBeFGQPIDjCj7AMGlG5qPQbo9bt/usCHMKiMmf8go1
ISM6nl6+xt36gqmwEymvlPoB4aiQEWSroYtSFEMTY/ILgIV3Z3PNLfOxzH4bCQIO
X3TTFpxprY5tEvbjs4TpYJ1pPF6NWED0EXXlhNz9yEYs7q44jAPl8MKrDHdwC6Bc
KEsaV2n+HzYsiijo5Hu9ixRfvJ0U3q6fwrvrY20o6yLfWlKIQZRGF4KSCtkSHoWP
4qC6txyC1rx5E42LKvQ2xd68wEg8pwk99d1kZcwsRrzKsM5nWh4PFNHljbNHlTo/
UADiunUlOW4TjPy3fiAhICo+eh/aEPZxPfHoHj5pgYYHWF+kuL+CtqndMF1W4pup
FMt8jFreBXCuF4tfdJoi5Lev0qxSvx3HEWyuzd1U2NEiWZ0NvBxyIMa7budnlpJ/
Yyx7dQ2ZszNNSX3/oxu1RJlXkrZe51QMHJroI1rFFyFr81/uX4qGMClPq+vCFGUx
ZGtGotZMhXZhYZjf3MJ6I4MuhA//sJLUqHfoLsfbCpl7qvarf+ckF87fHzHl/EuG
jrF/snieBDFeMKSfY2tX5EJFAxr6WJAn3ddSa9CDX87LJ7JPmHXsych+h8vaao5O
xs3+ECDBE0ueWkh7dvqQLeT4+6y4FCiVg9LZsfJSPxtDKt/AO4qlFjFRNrad4hvP
gJVMIWD0fVlfEF9M3BquOfzHpJ7Jpv1Lu3BOAkVkUFOQWptbfiPeSOPmI7F5mf8F
aaSfPTXGy+4ig/xMcXuQJURhAzyq5dRu3E3O9Mt6+s5Uz+IMukknh45n+sq0NCYx
LGaW+wFNSVLoYchvTo60pYMj2mSETtSN5XSQ4lVIOkDvs0dyn99o0T3n1MD9Y47X
5XAv1IJMrS4N8s97KkB66wWul7V2UZo1czwHNTo56kVu04i2vOVheCHPLFYCDT8h
peEGhBT0HzoRXNAje6+myOVPSbt5s36IXx2zb9QY3RUqoP9r2x4jTakDrXmvzff8
ngu2D4xz7saq11p1LjMqVbZ71YY4mRf6LczpenGfu4qA/Xvi+uARYuWBCPieCSuU
Vfabtp6Eq4844m/iqh4GsXDsHSzKgZA59oADSCjSStZnIe6M2Pa2DHP3rb+IF141
EZeWjaZvYgume0HecCHUO1cAyFGJeexde1IH5FgbkkRIdCnO8Vll95z+WTEV8zVE
UkoUmagKw5QMhdtBbXGm7XoIPFq7TfOkePQZVP+3wooZspP9q7cCh0Huq06VBQb3
rdde6IZ0lPb3MI9cvrND714W/WBhSufH6bEBOq9+VUfV5j9KJVoURWu+FSgZ5xjx
uYMJZ46Lz0DZgfNS1otR+YEas101WFl5Y/3sW/1dhTtDXnBM277tzeMu03qG9eik
b3YMp+UfQjUYYM31hmnatsdS1ghXkuxjtuE3GxdI7JIClbp6EX8yvKtcWjwTd2jE
Ep7hQ2MA/gR7x26swTAcUKzNEBaxSPVBGHCoPaoyELjiUiJk+FGN6GbLn5hvd8Aw
Kasvj4DK07lUwjpPJIhf9DTRSyY1nzphDYSlv2npqFuiZYIswg2EQue45DW+tlGu
OBHwZHmG8l+DAYItWuaeaCXvR4XlAldFg6oDdoD4mKD5WRrqeShHNTGXVojKU40J
sLONxccg7d5AtYxqMHiuVyK+ChxDM79NwB3phADvnikB0+J0yB4otKcI5H2vedeF
dpEObNCSfRb7bCVWl4oZ1qAOe8peciXE9gFcIF4dndCjFCk7uHq8NcEUA5F00q2d
zwUy3nz076v5bkcrutokuGOLjaAzLIB4hvUMGhxkzBwOoKVn+u5GIPlY1jY3+SOV
5me1+WAeyK0IXp1YxctAX23WVCYNBugQFrjnAFMR7s8kzT+PyyM5LH5/2jg2nqXt
hZydsf1+XqVUJnHtCGGZskV/H6EonMIn8EfwS5AXnXTeBMHqdthJ8QpGv9zuA0TV
1VSQ9oAF4Sd27Cid/rU9SH4Mhcit5GGsQMeF7+5peNve3ers50YERMhQMQG1HcRm
dUoYVATNhwtaoD7Uj0YEXH3orsM42Rrtc97GM2Cfl8tZ3XLUEHSbH4F1FFvnh8O0
VfuzlwavNyVloFnC+TPm5fXkBeUckUS7A9cpCw/KIvEoVdHxZWlMtBoHlsUSt+r5
zvovHEZowmK0Y8Ons9gGMrM5YkUW+5bj3gQU5eOrk3wlaUpfZCeghGQ4weB4p+KZ
oUpFJITrgKO2i8yTmCODNu/dGO+cPsZkqUA6L/YA2VeX0PSbOXTP2uxat/YXooiQ
TBACj+QOZdhWPU7el8vKJzoUkNGSzX6qECnWctOIsPpjyuYPA4DQyZvlLZUBKscN
Oa1czJ3XzgTWnhXEipJ/M2rJ70ARx9e3WeEmxfuhXIPZvomLrPGhtLM6AjTQ/HC4
kUWI8Ag7IgqRskcemEvQvEM8vuo+/EYUdk7TPGK8LH5dbbIA3dCScLaY2IMsIZhW
j3jxDbiPKo4Sdgjx256SXUvLvtasLJYX2S7cqDZrLTn5TAu1Wo7gmItK2St8W4Z5
lk7waPfj308KLB7wAWpL5Bs7+LkylwOW2z8ioFtQIfnRSPhTPWNEJtH7U6EPcQY2
r4EuSAJ0WDJAWtIGJupPPnar+CmxATSOVrL5ScXBG9zjWgacmnVYfU1oW/5IuLE1
MX+/yS3jYqB8RwPoc2vFMt8wNlBA80b1J+kHbXLs3rcuqkltf3AhGdWZlCmuom+h
DF+kQ36AwrATuFRRrLdXOuGmPI08EhAH4+mgzc/BWAPKa+o2zd+pW2vnCOg/Kdas
Rwhsl68MQqukpmiqic/1ZZoVcZA23tKczVPQJ5x8H/gY0dKS5Gpvsdm7sgdeDZEb
m0q2PfEO6nXhyVQlC3+bjCoorUo4tyubaGA7QFWkY0oWS+jS3dXgsWf+/47NNeZX
Kok/3lKtRx/fw/Yl5FP++plNuh4d8i/e0g3LrSiaU2g4iSJhSNwdznylhVFBKikF
Z7LTC4CYZllYAt2Kr2mRBHbfzH6T/WwJcf6dV3qb6ydFCNakCplpt8drpQdcX11y
bl5zBZ/0TIKnWzhVrBW7qCZiEuB+K7LaBa0+sd310Sdv2RofL/fGhNq+aN+45O5y
8Lr9BOCpSNrGuTp+1xsNh23pjyPgIeBogR1iVqxjC2VpswNHoUxD8XLB72qiJrK3
Yqt9iXAec2Y8olUTzMus6Lmmb0V+RA3OwVXRzbIL4CKWVin63lR9/p6q6vfPguU8
QXXOIS0U+H/5VcsiyQa8GLxyWnxe2NnXOpSAGGVXs+7zZPLsnkZ80GAFd6lSN2nD
YvcPnmmeaX7BvSy42ydLWnSzqoCwXJWL9UdE2wNbV508UVbsmEjK23HJ8ISB8NLf
BPfqxlywJdFw7PoLEbZ9I1oRMHyVqGG/CEpKnU1u4elMiZ+PtIVRCIin7Ja9jCt9
NAUGlvPwBMVKF/claqTtHc1adonJp3UlEueEdonBoDkLHKvXQrJ5RkCdcWz8zhxt
luo7DTpQ391qS46HDgDGPuaSbF7smEmxYjq82LByALxUBFS1iB60nXqgypNXAzNl
4qKOTQd92L8kBJbLLeKMJBUHTF3X1vngEiaeggd1jDe1HxhGuLnpm6L8PQkw+fBg
9Q1Ye/m5hbxgCdx3UVdmz5ZKE/wLjz5wF8Pu9aZnaECHFWiWIyQhQo/pg0mq3FGG
Q3EaMEfmy1+v+VRs6NajVrZVxn64jZ+uNl0521/YE5p4wTxfIZoW/LF1HQ5O8EtV
OoDlJck9Pr2pKbMdVGphOQjMWFrrdUQgDG9PMXY9yG48ZNUmCsRY2ncTz+l7nW5t
HVzR2JJCr130Gfj6rhGa+yO28VD2bqzqE7K7GRrTjuMgbrksdObcZKEeCFrISPbd
VlzbGqlqHJkZcOG1SQyN6FHMjxLKJuKhTd+bspNwNtygKivUBmaN93VwsT9TWP2R
v9mGbT8YIHdNP/4nxoVaZAUkmQHuM346kjL5uFQ/Ug+EjM9dO1Zh686GqzZVsb9v
FTBy6Be3uKJHqGh0f2QfVrPEKTslazI31IMX1kjJa98E6zPWzYhqaEXfeN0fBhne
wNfnh4Ddu8V0rLK/jumMsbFslIz/UY59/UoBKCQ1zzTD1F92QA3F+4hgXTO3HDKN
zIaJ9NSasg0ubOINXltNZhk+i9J1g/LyKnJ2ljIALTXc1yUNQXL3nY4Tm8pCd/3D
IlT3Hgt1Ft/uyV+DxPJV04OGyz/NspxVZWHN74rjZzUzInDBEwmNSH6aS+1k0Z9c
9JJZKkubMV4esQ3Wq3pOFjj3LkekOL6NC8WW+2mWfVHtzEiv/6wGlc1r4o/Rm9GQ
4G90dxtdYyw8hbRDO8w3t8iVauR1az/w/v+PdmdDJbSdjrJuBrfB/rFz2cwh/jcY
mqzq9LYxnqVltggTbnHGKMcBJ1ubyl1Fqq6bfYOjDjEldRLf36UfEgsN9M/3ydVy
mgkCu66LYEhHam3Y4twXUAl4lN4IcT8YHdwVcFJ3DVXS9lbXNUC5ujedxMMK4eNY
gb4OOcc9y2iVnBbeFzYg6y81qkyzPf71QMUGaJLaodkLRKMeGd1N03QASs1bDu0W
bVJVM6DLpV48qNym/ofrhvD0gBYawwEutIWpB7VzBwuk46oXLY1uBWLERNHtxpzL
XgD7dkhd2KxEmI1Felvjx116cV7p/UH/sVsq+rDBqClAybFUCK2fOKO9qM0B0oZc
zL903KovzUKhkf1ZYdUQ/NLHHNoTSHLH3uzRtAS5vRMw55WVFs7sduRa+jVo8LG7
f0OcVZAguInv/i7odGLd0LgOZ81yqM9J2i4Je09u2aWhvD5O06CMoeTd/yIiRTCP
jUArsCWrow4wuDfSEpr0QKXPM+0oq+EzMItGMVkIxeZh7BVl3m9Y8e1ke8BznIcw
VpTTGO1iL0GusWZtzwVF6AXwb18lBeIvSoAziIn7QqJP8Se0TUrBeBHdNvBJPiP5
QS5vgahcIWY384V3cstKeSY5W4/99E3t4nBQqotO+qHwHSFoNmkoCV6qPzoXEoIt
Xhs09+5YRI9WkJS2wpSFGjHEDzr4hbaZzA3j2X+s+N7DOFvMUoZpIjVGBiIm9PmV
20KdgJQn0KB1qHFyqAIgVaBYY0Hv6jOEarv01k3gW+KYmSAKTFH4B+WUE37hY5MM
EZvg9J0iTVHY5NEQS0eeYZR5l60s/mKMHv8c1oJ+K7B2pJWmuu42GTno5bTriFIG
vC4d7gJBB9kvqe7y5mlCLIkV0WKtKNXbPaBQti3CRCO6tKyD6qOAR1/dLBHYznWr
lGdCODhxGswvL+qsPUwtmfUWqkiMJdRdLEDw8v7b9WktidkvW6IpNappfKRULou0
gDKdJMnDNp/o4pUf88LlCW9Y3qiMPgsrlAR1nsThsyGoCIN4oUGIM0+YdNsBz9pz
b27SFA65R2zDitugDW0IU31aC31k1zkhBN6QqSRPTxoLiGHYqPeJZT5KTh64hBaY
hm5V71ARZy6Etrv0WMVBOtOdsTHYZVhXBC7boCdn+NzwrLg5VxXcoAE0liPSQ9+E
f97/OawN8fN7Ix4chu2NgNRvmjlldAOasbC3ZlE+rEk3iiKePGZjgyKa1bwygNuq
ykPl3+ue3M4ECTyOnYNHohAGkGRjtejDR3LNDr2422cVK1UF9+ylOQC2ayaS9Y6U
EzG9HevvMlCoKtAVb3hOLRK/9uzgnsk2sCpu3p5bQwGwSkcpxc+if/sgksJZ03X/
xxRd/hOjEvrkFhJ0W9ojbeB9aLNwjTJ+AsSbtvsccFW47Oy49S7gs7xpEH81DO4T
Pi2UW7ondyOGsCdLZsBNVzgRmusQG4QiAOEXsERy7tHlADoZw5h66AO1NRqy22N0
e6ndYzHNEB7zjAKdRK2gxvWEAiDNkQqT7F8b5USN4z9Rn8h3g98t5DYIXSZQ5Ufn
uYsCTDGVO8TA/JorxtH+taw7Cm4jFDqoW4RH1nuSAmmG/rw2nAbflkHDnWQ555rI
GumcUw+V2AzfskOgm0o3DxnPEbLRTLwkupcTVJE1kYnJZUiESCh5HonmxYQOQS4L
LGyBTDEAdclS6grRz6SylLGqGUs+dQlYcyJmRIVYvDwQeu8T2AI+oASj8sejoyUt
mI3TyxLHxuM4uR2fOiQkRLc5dg62eT+DwDSod25morNNu/ybXlmaKanaM6vkTih/
ptMcq8FKOh72pc7w3SqBj8ILcE0FH9XydxH0Cc5ColQN3AQEU73CqjL9+j/+7SwX
a/VTfBd333LB7Yan5L3GKL9JUqaN49DPT2KBtYQ0mr6G8G4aOyE/0QcNanhO/FhL
aRrnBPGy9u9/t/eB7jm2/NY1kMJTdfU5wZUnP7W0y8WF+Y+EDFazUHRbPby0IBFI
0k7t2TSK0eFf9doLDP1L4Hy5YdzcRvnEmsBvzywOUmCMLwswgJLGfYyVuQb11Wrj
OgUSdCcx+MfCCYicOUUbhZ+r/4+i2ux+TPTzbRZQTrRsYc9WOoSVAIxVKLH9+ZfB
/fkiJVZ0S7MQ/T7BlzS8hmX8oTbFBTfMcCtm1LKv7WfupEKM0I1kahlCiprI7tXk
wNWJL5hXwcN/AlB+eiqNgRF6ZN9l6x2d1ecfgOV4UhO9itkZ7VlCq1G8brQiDmJT
oifm7/l+9coUT/FnvDTPUH4Em/XrzB31t7LqSp0FcbW+muhtMxqFQVxw2SBgP1Zm
2fnCQ8OiRtUhCK6UE7znmNgdZX1pLUDryRxjw/hh4X+mWWqufavuz3LFzC8EFN23
jKtIk7G3EnGLCfpDzAM7bxxNdWkThZZRPoRjdWfMwI2z5fZOoM/naakXP7cyxnh2
FCkvDUcHv4rFR7dwmwc2W2yNdjT0PptNW1+Hm4Vm7WT9WBtUcCkhsuLzKAYCo3WE
9s7yN5mvK7WxmRj7sZ04V3bvR7/PLfm+0Bnowl0QSdBL9NGHVMoUuvAOGDi1MziD
I/MXB0KkEJt1YZJEztI/6q5/s2frfjOZyFGrouSwtfGKUyE/63zFhVRKhgrtuofX
mN3IS4r7HgojgEnZn425eLzhb9gF+zwrLSk1DdsOIlpH55fTa1HeqybyOLNPq2FB
4yTxyD3EQHKj/7AB5YTBUBx+XoVfsGiwiK3q8qxQVFUDHE1zaXOuMhIqhGzK1OHP
+oj+8ucX3qIenV6lvcC6VWP1rrLKUajWjd14V24HrHsdZFhglVF9vVGmuLOavc3L
HLQPrLOvWW8QnJEgY0yP5Nz/j0A2KkX7LQKS+u3DptaraYysmFL6Cr5BbWWCEb/A
J7xVy/nogSAk8zysxrYapsWh2aFGC9sterMNO1469knJyBsSXm76bWLSpvln9E6o
zUyh9JhBBSmr88L115+dLRaTV0z4dMnsORBYyXReuDlV8YsN2RECClBDwg8pBYye
cUcM9L+l6Mr0crK078IeiNjuDxJ4y0ApeN8Vp/3+ussqSoBh3cR3F96vcYU8j+YS
LMRgFzcxF4yAvqWPH0e/AhnXh9DfTCh3Oty3PxzC1gl+ECSWyGO7ZRNbMlnrYuhg
F4HXmLoOGdFDOfu6rhg6R/22hogpoqhFGV/YMkpJBIMg8cVe/flkb8GH/0+dmY7F
D2skoe9NkdK6wRxCfAp4USsTXzq52Fopgm4TPklkIoTsCqc02cEU2je+JORFBwID
vRFeNhAJfb7Vj0oIONOnztPJcb8T5S1PClVjeO4epEc/BtjVf1zGhL+0MWoPC4AQ
X8+PZnczxr0xLgw77F4ywO0wBKE56a0bGcsS9H0YzRJmmsYIWA5gEBDMvOPZp5Ot
qxsnAL5XusS9JJ5CoXLQVMIcTYDIkx+UWBqu8ZvmUKHAk9zFQEnsUzQUNSIsKHph
48fgkpOS2d1PhkIhdvRpGD4baj5U0+PcDmNI6HE3GzJ61GW31B0hivKXb0QIekEE
EfJjQlzQuJx8JGvqlmFTw22HeB6QmSSEJfHEKo5n2qkSedZQ4QjFgX/Lf42NedZi
a5QDpO/48DJDHpViGzNnpNsejZPn0DaIxsEM1bzO1Io5fYo9ISrBG6Q0zIwX4CZR
4O5AE5Z+XRexvX+75VOrUxJVwmkP5FsLU8R0fbiK0cDupY5Q0zVyAkTIvRU1pi/C
flklVVXl+GALp5Ss49V2S0JKX2AlW1p8XgSlFBiTjuqzk9dXho+KTNk8Tzrbl1n4
Ak+bL1lCUQX+08xQ6J2byFV6LhSaHzJVG7xsQUo6B5waGGCTW1LLkoYmJjCA9c1B
avMNzUOlmJDGUfqWEb5HD58ns7IX9lIcTh/+1wYJ5aZDDC+aOzmPDtJ/DpmQ51bq
jYLstQd4EOXnXOVrkmDa0l66sQitDuEwdtFQV30NgCaWoCmdS6a/mCIbWgFcGcDd
TI5BoqNDkb0u9HwzZsjvw9/ykw/CB+9iSvHx8zONi6JZCzarrV2HyqYj85m8Th0U
vbahh58sCfIKdzUSEgWh04oBdtSpUVD8ovgbUFHAXIOgW6xP0odPXZIpm3xM4YLj
gf17cUvEeTe661LOjUYK8qKPB6P6+AGcU/LFZbLbrNCEp+fv2JoNoFcC0DCHhJ1j
XXaxI9p6rt+qOThNbCO4z7y5rMh/MSQ0UOOK2G26nbzsXB2GmOyxatKxDzhJYmdX
o1INgWS+2c8c5ulgijHXpIdun1FgJ5Vch2AjqCz6XPdanneKSlZFo8iWdkSNUSbp
OvEJjGoevX5rpxTBc8peUc+pVhtPf3jaXqZCWhsQ6Sl/NOirHkz4+ezdskBp8bvJ
3OSuOi6KE2N4V6l0UhT1YjLyBPDBRXWKlHpU9GTPZNBq0KPjRRTzFGsRyg8yh563
VNQQUelrKBfLR23Bms8zb1QuV5GQOIyCpYKrTeC+h539G2oskmGoNyu4Vt3pVqJL
DD2mAPeh2odgy7HSCxcBY2rqF/Scfj/WICRgfYWVbWhWNQQ1zH9LnrQcXT/OfhoJ
Ab3U+A00Oroxp5W1irDr20vyjmojghuPDuSProf7CicU/ypfylHeH7c0hO9bHeck
GU6a6EqUgyM6mLuNxlwMIwzMw3iDGI8s2vjFrbzGFoFlpibquEiV/BoZvFurgfa5
pPKgpMHAHKLxMsS4Zckzqid3yWpOIit+aU6XIzE1M70UFbuhYuMU4OziA5EZ/c6A
EKFN2lxFu957quGllrlj9A+P0imiyGfpjwoxC3TsRrik6VpIZaF0fN6p/rbBdRrg
u3tk6N5tePg42jyN+u2KDV9F+YkF+6j7VSrxGqUNrxL8dEKIv15OEicJ32OsmxXS
BiFzxcmWps2JFEUi46RGSc0ZyV6Vr4Wjo43Cq9hdvFauFkKJ7sQQA0cGFmBpVz1Q
Jlas8BM57ehwaFRwDM0u23HueGWxqq8Ah0sc20kBCLOPC4bNqK5wsCOjYECeqcwp
/LxwmBLIulZoNhwdpEgp23bSDLbo3fTdcLnQYPRBRqdeKm82nHIlV2Tbpyh564ki
AKkNTCbVec8qooRjuMRVqhEa9vXALskhYIUJDxBc8wgDe9/fttqsdHmKCUuT53CK
BT+fEhommpZ9z+H9gLgMvyg4YSS9f8BNla+WXq7OsCqZSdofn4HAaDRuEM7RKGec
3n1stfPXtDFqnsa6CoJUwxb5JAT0BZ5d5etXh0f6bOskmthFbXv5e/ls8NeblbdA
pHDhg8qlfbJRzjsyBXYmWCc1NbKIMxU0eQGUq9JSroBH5qij4p7lkQ0rgUYOHNfq
IpHWDrOkGffY/XXYIROv6ivFKKYbG0MGsjKZ5U8grwukBGR3tnmtfBTWP7NNGTaJ
upUajZyGmta1bKOfMcrYS7iFdWfx3SyZcy6i7nJeOwdAwH3ZWAuEIHc1sqHqK1X9
ITQTgu1fW6SaTAc6LbkVJ+DTo7+sL71fqsPtyiVqJPPAzuSWQi4FcPqUKBDSlerx
HO6NUoTFl7GXbsGQonRiweir6ipvX57mb1bBF1hEFCCVIGcGFv83j7vrsimJPmHC
v6rB5slr3yUYmi+cP+c4oTwRz4V0R4N2LCzlyvSpRRk1gHM9iES4GLytGl1WjGkH
O9oFchR8qPnXpdzVNcDx3sE69DdgTgD14rHyf7HDxKDZjUvX0sgTSgxfn4ZtFhBd
hboBM4i+CaJVjn9c1pGG0uxQP7jAqICHO/WnD9FqJ77KEJUADY1v1lUmyWk6ELId
Wb/DmZW64FpzTQcNy9teqIgOWPRPx7PyPoX68ykG8AMrCWOQpsuJ8oOg3LTj2n8S
+HGkoNawLFq/ggZ5Em/Tk1oDjorTugO1N7v45VJWa08hn9V3OyjehwE7duKKtV5W
/MnkSwLVEZbHLnx/JGAP/SaiWvGbG5X3RcWYMMm5u5j4G35ssZau78DsjacXbGSz
ovL23eOvxn+YElLvg5oIZ5w2aTc4OpejDf4Srf5mEw1XIiUdBzi5JFkQI4t4VDL+
z/fDBGpWBjLEUAEejZrxhD2BGvSxr8fii+t8kprqGUAklJdSQOIb4/+ug40PpjFl
iWtrvYEjlaVQz2oasJvjH989AUokCR1Peuk6dtul++hoa60J/uCmCQLBvAiL59EF
Ou/ESxBHwcUgLH23ONuyWUrymRRQdEajm5DcRpVozxCidn/yKGKfiJgJEV2KleZh
Pwhq7Y4a5mpS2wpdTkp2RbL7trrpLspG0D8a2ruCKUHljkCBBulLccNUiA25Pe9w
XcRoEroR9uVPnv71GnH1mxOnkG/HHQzCN7gcEs3UTb+nEBoTGjvoNv2wZ4EQi5En
FIY7nZg6/joyEl4mUhpHoisNEmVjYTd931e+w5GVDRntFYmDSIlncWRXF72je2tF
SQ/1qr+neq2heSDrm/x1w6SYkMktopbYnluiEtp2KRP1+pTVnGikMowgVPLslOBb
Br27UDgrwJURhwIonFcAuZhrV+c+NIoL2Bi/eMmKwT7JtW2azrgc8U8pehu1YPx6
rdP55uDZwC2gp8NbL6dSD+/vPHbmWE48vgwvB1xXr7VtTwRNC+MROqUs8+WT9ShT
iE9BjEqH3EeRqe9e3qkyu7dAJWxGXmiSbZ6EmhhM6qph6cGreTz/hYg7YRuVqkDy
yczSyyBiLFwkFZjB+9rAf4d4YGX4IBIDnQC6SFrawvUujwDGKlaXEwuCDt5p21Oz
BrEr55jJw/VJvecQVj2biYnoktOUfohNReIgVdMHRwajmy7xAK0ui8GnLIVUyMwj
JQTNcU8VSRASoJ2KaSiA4lHdLLT9uVN275HdhP/VpF4HJo48pzw9nwDv5vUJeXVG
+F9g37gyFua0Dtft09TeAXj7J/1eGCM7GcRiyQzsHQI/9QoB00Jjkte+NejaSRNZ
FwNNc2AaYieyyDC1e+bT6vTHodwTMJ6y7zXFMVj+w3R1TlXm6MupHtbain491UP0
K4S5I7x1mgpR7B+D5K9d6VVZnZsrVm4stEX3hqZIwW0+FcArtajfW/fbjQw/9M/x
ney/VABXxhoa72sNxKPLLCYqpEsX31rTj7MQwihG6MqQN/Ju2QobyA1pDIMUvR/m
abFH/Nk1KLIZXFlzYIS3tUDB1RIFUqCH5MRuJXgHZEdUG1BjTYkP44Qlj4/FZJu5
wHtx2qv6uqM58d97XkgiqmPJcKt/fEqsdz3ZoqB69VIhgFP/qPv2ISZ6w4msHL+q
TpgqSMWZZyEiQrJrAz4iSaWLNwOayEfL/iOfMHfhgFDCDM0yHjpKnAD58toxuJ93
eXKbD0N3RnoKDz1LV2o1eOAMiWgRwJQrMLlLhvfBTMNsn4cwS7ZNqY0YyK+KcBqJ
d2Tc/QJgxGAwiOuYn0uLoHclpzvIbYUNLBkoftbnvEj9q/WPD/hpP1QhTIrVPBBA
g7s20moQVOYs9/0zblaJEi9Si/qupFyEEiPYDfm1BIWHLrwZFwJ4kkagk557goi3
WtCgahTqKg5yhot3zTfK7dswsZgzZS0EjbF9UNG8ooysdEEP+r25znP9Om9tTR3Q
4kR8oHBTbMRxJUERlbnfu46JYDn3ZvE4PeWybjD3VE01VSczaWwXwhsMctzcJhUb
UkEK609RB2JV6IWOxq9sjopfVqHBQBOhFoB7cGxLqJuD4p4beb5VXmvEmMs/abGY
TQ3Vmmw2ybXY+WvdYlg7QndxHBnDKs/bzpfw218yyYgqVcb9vO+bORXgNaPq/IZb
e6aSfijdSkqfQpNxJkXbm/2AdXgnGCX3zFvJxOCZPjIM3RZYnHRws/UlXubX3zZv
yaCvWyxGbwOYWQw/h7q5+zOL0F65H5kxleGMkjc+8jilz0RuhQUV6v6APTZavw6h
65/GEsDMtv3OJC0+DSg/r3YUuMslVGwKiHMTiRf718pB/I+hV8gk0n5DiL3WCDli
AHRiXypVfgM+a5gLGHaj88slHi8MzSfvb5RDqjqATquO8mGqV78YrsNZ+gSEzG0m
uRigUOuPi1mkls9B3e6tq+OwVyb3+asxbKHhZJCHUzSheVNfu4hdPc9g9hu0hApA
8Ki8XI6JnWQFuC25YHjodC7IM1M8HsLp6/23oN6UqLoOlo6lwbheQ5HYZrCus3jI
mDl32shnnakX1r3l/JGsGUHxrvcv7geHBa282E0Fu+RqG5nAs5pErnwdE2DGijqc
JYjOYMbfZGRAi0Qugf62cM9Bm3BcddqZVyKqb0wp32d882TwatBm+ttBQwpBRRI+
AXNiXC3GM3Yn3sKcbvY6YU/alsZYDn5WJQuKNhFZT1apvWs3diMmtuzxj0Hhy0tZ
01T7rhDJWWPWC/wCRAdA1Z8Z0t8slKHc4Qa79CcbaW0BpmxFOmGcrLbfixxOis80
dWKjDSShrBtnBwBqnXErAFb5DmNfN3jOoVgIE/3vXth/Go/dsFp5orKr5+LNpk0I
GHrt00zK3ah9waypMzAIkXIDx25kmeNcjQux+zSlD2gCRsdY0+8bYjAc7XYOqjQM
BYsFLAh4eR0foC0kwc2adss+4j3B0ibX1exMF07mUmJrF6GqhLCeyNFHX/awJDvG
pzN5W/zhUGRfW2ne0hn8x0SA8mxFiH0FUOkJ4d1Kl18xGfATmS85PhB+daEgq+ks
y1yPTYCR9TCz0CsnXM+6TWLD1f5giqFT20KuETR5DMZqHFCXxpBygpMivr/yCy5m
1+YSVEliuG5dsOeV0LS6/OAlTOsMhBif+fSI+LlK2d1GKPXP5PwP1pP/sHoqxaxX
HxypFqyqIKUmflKudycu1M4oUnIW+llzE1p42iCn4lKtgS8Fdj+rIqDUsGrWZK8n
4uWS/KdloGvBvzP5Zsj2shLC+qaYhw/eLRf+87TXRVFh3okyl2E41SHzsTnZBLMg
X+y9WomONv0YoVpUsE84xYaeiChiDTKerNpNB9otPbnTQ06XYlluQ5pB+LnrFIUT
oOzo+EM42Z70wIOl336QYsNfOoECAHvpyifb8PB6da5Z70Z10oLsJ8JZtsgi/AnK
CdijoU/Qyv0Jt7owXvUvAUl89UhloHmAyUGcPNB76jYdRS+XlU5gpoddR5rxAn9/
EFxtMx4ZARCH0+M3zbPwPoI1VfOcsp5Zr8HXrKc69QidcI9/jJj5i01AdmfBdzex
ZvwGJMi+/YMnFRMHFfrsIjN9F6b8PQ26bOy5tjnUC+8tAwk0naOXEWERm/n8fKVM
MThcfiz4Y+yCjn7iki2tyDK3W5BpKzZLbcCQE9c9ibULmE6znNOM5/5skigegXYS
opd95YX/3oC6UlKRGyY4ADjjVqXJJGrnZ7p7RB5RSduq0olOLjmrSCs1KwHdrEn9
8gCrlnLGhx67aIPntVkf6vtq4HD4XOKBABFhyPyh3P13vpOAlr8qKcw23SlLwLj0
XTfk/S+/yFK1QIRo7lquvwQpD/l0kS8+6It3as1tQALfhjLzIQKx6JAp+lBtcsDy
eR/SMhjLKWuid6Ea0im10riBTsirhSOvnTVBtVYIoWbta1yZrowtm9hyOXOuGJZ8
zYH0+Cwbekc7n6PAZLq306MnRdM2rnJjfJt+nzG7WNTXtFJULg5EQLS8fgRwh2Oa
QEgi3NN3l/Kuk9SmNchoGw4Bq4GkZNO7wP4MSsr3OtItx0/nfEU9+v0lOQIatAFG
VULqYPBF7Xp5R2CQBa72IgzA7IVbKukrnjZfqJfLPXxeZI69EfltGWocbQKxZCPl
qA+ds7xHeOZ2NIFX3Vf0h3CyOrPn1AyS6FvXeHg/AH88ByZcACGye72usQowwDNE
m7xbkUYKydiAyn+ge446TkCS1NKSCXVULMO9ADJLSU5OLKwf5K1JRp0/JgP8ELax
hlE3RMjXQs2YzHl+2emkLxKbdw5fYXq6QE723RJzIHFkuq44ExOn74wxOXeI/LDv
pHvFKdIQPyx/f9aQ2Vh4YZdmxlqVqezrapY/VIZDuhThS4OYcWPFMIKojgBXURzK
OkZ+OfDxFA8vnFlxJ9JMWwzQjXJjePwIjuxYUaetmwPkUbygviH1jVLI+CO6zuNL
Ci8bOmBlM3Xs6mR7g+/w7er3hTsV5GV8s/H1S4uJjDVAuIqfkejt0c+wQIrOw4cE
Lxb+v2w08CawwMBcFxIPjLF9SYeRiEL7S1aYmxN/QicWFpySkSlMtxzdNyis453O
gWYvyeGCyx9oHhFT1adgAS5zdNRfe096J3OcZ14xT+e+OUuJYLn+uXyZXfsvXUF3
/gh6FbcnhZbDhv1v6+G7J+e0r5wP2nITbs5BLzNjVGuH9CKUGEE6CTReLFsBMjz1
3XyOFZx/yn0EIVrcJ1PjT8aL5w5pjksTDVApuLtqQtWcKXDK2+f8x3ohZ2IyS9Hn
uTMwdDdx76wklFWrccqkmS5omPHl6H2Ous1e5fHuFUSfH620BEXtxksHZuBHpXHF
MCYZQV3navastaEG0BzeVwaAxjqnNVkgNdl3Td/TV5cZNMODPq64QkduVlPu7pca
N0HhhuEHzfK5VkBIagCPL897EwASZIOJTcDwnZuB8Ms2+472xplsj6OQGVfrhz1x
twsC6ALLdQZ+95Obli+4Ir+XSgLXrNjxOEqJUZfyJS3zQwqayoZNwElac1Ly3AP1
GePKkuCugtBZz1CqYkAH+EAVbPSWdztIvlhFpj2PC4N5KrqHRAcNMCwQoLA9JiRx
ngnNeC82RHS4DT4OWbUrWLUFpXnubcbS8vO9fYb2ZCMcywv2OpeqpVY3UsE3UrxU
bWp3qKNiqaXX/YpAVtAU+3PEGG80VfBIZtkdZSTtEqQBJZ6jSuyMSqeNqByYCTDY
MN2dNXql9nC5kBDHoYbhA9j6XklFRzSvVdp12/G8z082tifc3EXY9SJ4325bufZv
krpo9YeAZDrJgVDA14EJH++3Qdej20B0GFuOYrkGifYzWU13+x5qrvS4vvYkSpRA
1/Jw6t+YWsGNpz0AJ2P7gpefPKYWS25vhNyVRaqa7sqLt+0x8y9EnfQisZ6ZuIHh
/yVuxvrThuU113agT6+xJN7LIE2VJ8+Qe+LFkNPMPBHTCobGg0Y1geXTsPs3DcC5
8lcnp3LRaP7Z/ks2X03Gvf8Crt87WPSFqt5ErMLNcL7PfDStG6gew/EvmMqHPqGu
lj+PxizCc5FyN8d0Iu2MbtPKLLEf8MWTHdJbRL9XCordt0568k9xtOSFruqfSEOW
BfhbBIqLMopMrMYTOKdBozpWLFdnsYv/HlGF+mcCXKQ/C2f8tNG9o5k3yTmb91iW
Aj9ZjYoWuslnSQ/DGGTmN1nenvhhxe5vR8+3/pXLqWgogxcvp6YZScqr1SgSvB96
0VUPdn8WqF7tl4DSlU8DqH0D3xFiDR7KHb4JHpExX5/z6aZMj+mn66rEXuPG3Ah8
hWb7SEUs7jUecUxNnvZdgvfi4Mx3hJ206r6HeRAI2a9CRdbAd7QYcu4I35TsjDue
RhC9mD9B9nWsqwhZcJ3MprCUvJo1UnJ9Bdmbj741N4Bz1PLlxomnS4TFJGYWwx7N
VY/qwhRI1EAHfXaWV4NMr32JPzEETO7c2+JG0o5xMnveYsWlYqQZFXxUoVETOGc6
5kktUcQY89Bm+A5DbvMVLCd2C4opLKc8rwEMbOmrm7dpAmD5y5qcgr9Rvn3pLlPK
6ZzKUF+gBWwytk8/FTuGeoYmJo5lk+3ZvahLK5aqA1i3WS4NIPekyZJVruh/IthO
KRk9xTK47aa2d2Y92Im6liIByCGFky6yYuZVRNiR1JyttZk4YP7Wvs0A2WCjJ/sD
Trln1Yy1RFo9msCmeldt1ziHmrs16KWS/7v8SPXnu5doAF8B/zvx60Arp3YUeKTi
s1XMSgg3Ak6st+SbCL+AsyHuD5np23KZBSualJ4Km21bU3sGbU47TbZDfV1sfrJR
FQhLw2eigxF6blHU51cvR5PFjaUN2muvxpKhoh2lBLkDF/LBhqWeHiG/ck/gWZfm
dlmGIQ9KMUgEiT7ttCH5H3fNQGV3hLzDz+wUBTmCsjLhPGVbAoDFQ2Rn4IDauCTn
Qsi32Eqym+akuLpuMeAiPR7QtqC7rmR1lTF0Ces0pWUQ+le26m1kx40I7X2IpdEe
QOcEyML3yEFv7+or2ynEmXf1daR3jr98+d9yMep0dK0ab5sZAVI/XsnLq7QtYsv2
XKX/cAvw26V/j9HUngw5TgVd2FQ5ThBeOhUxSq1Hr7mVgQ8KLOGuRI+sD3n/EcS4
1Xy9RtsCwijBwK9erZDBQBJZYZ5Y8t/lQmqYS6cIwvMnI3AoNL5vYa7N36g1bze/
HZH8dGbL4mpA7MkSmVotQ+IQdV3LXqm5upqjAdvxbrNrs8PTfRaSO4Ecfu4xrK4o
ZKN4TTmrYxoanQK2/4K0ms2Dj07Xg7XuMKwj6mkKtMoAuu+6aq32IPgmwq7/emuP
Cs1pToRboHmaU+KwDsuZUzNISKEjMmSahLlOwo+/YhppfvJIYblFFBmBvh2TMxlU
77qXbj/t0+DOfNRCqmXmp9EcBNwcN+1YuNf9RM3KHis50S33ePs08Q4t6h5sK8Ec
4tJY9JVPsq/sQp8tJt+rR/Z2fG3N2JPsZonilIkEo+7gXYPOwGwWsZvf/M03Z/bh
X8mR/WJAVuuK+b1cYZCQOe9Em6KHc8UBx8iFVkXLw3ARCVRz6dZTGtC3YD8cDtEY
RiWBgY+18+dRLe+nuqP/ZWJEzh0VomeR17Pu4ZYxMz+0kTVeFoJ3FJI5tekQ7uVX
UorEAwvko+UoP07SkJq/LJ0tP9gEhQD+cE0qfb6aDCcFBROLJyUZu1JgmSo50qvC
ueipDlWszSP/p7a04dBRRX5/pBeOMIRQyVWMqtSad7YRYrLIpjpngUujSofC84JS
X2Ir0jglslpvkmVhgBI5MoACU1gNitn9UsdkXLcOZgtUB03yC3EvgEH20hG24988
vNEfxSlHYLTz6BACB4CbFYtioQiMt5lOxtmaoBp9ibXtcVw/aVnHqAyVBveUPp42
5nb78c4kRKc9rv+xLsz5jy9LQKwoB0I8UXHBQy4EanxLPVZqvHwbYlPA7hcM2dPj
ZcIJhDecsToU5iT0oN44PsulBRDnBWSDa5uKQE4EHAZK1YnMXodACvXhC1e54UYZ
E2oExxGbIY0DU9j+ZRKicogFIaerY6IQSgIt8c0XGnOe+17w3fLmxSnIuhV9bNPJ
SrswxnxYADU2O3dzQVaE1I6s0AQ+9a77N5+RrdVhQxyYhDlbGd4bpQl4j+5oga78
YPVQyOZgrGBtU+UBcW3H4ebDY4mN0hfp0tjSOLV6wLzg3VJconSxD8+qH4+EnURj
j2FZSE0ydZVEWV5wX6dk8cQZBsasNbd0ym39t9wfolQNeykM0js4Hw890RhMW9y6
Cm5ELD9B6Nj+LTPfeyY3p8XISxx+yvUzCriwbyic3CmYzh2vw1VhWlEV27gfGw08
zKGiOImjv2Ihs3rgjgNrowntJF5YpraNt+nZNcUuPLo6G1dSFYNVWJHGr7Ebi+3I
rHvpl964stbjcP+8u8D2sed9AQUO4LIzl2JNOIlM8EMQi5vrt/wOOHRuGUKzEmK5
avqBVF6X0VTblh8D4Yi9fyhRGXtGRkaaijxCUpBhZXL8e3SiTv2mBSWGRFjhotVA
mrGwUGg7oXBAJ4okXiqjJC5thuh5xh7MknNlabqGTtkYPBU1PW2M9dkRh+206bBZ
8WeVr+S+ASIbkTPcQ18XE5iY+8f3GWQ2hZV2G4WwpssWy6njHP4OpFAR5JuD8JqE
bILHN1ovNqXQylHyK43vxFxTuOAAiVs8dWjRyqDXHW3wEk58p0j3IFqSks21wOyN
356JaVH4KHc8EuKfJ/15Axv3GwFTEt7VHl5LatRu7QPtt8rXLxKGKgCJMVohmRFS
QkwSFtccpIoxeS6r1pm4A2z/tXy43mNyPUt4KGtaAZb+JC+U1sv4pRBlOj4Oredc
GzXzYn5V19uAWGQAIk3BsejweYLtCfdzjinJSlNP+eHqkjs0jFSVgvZCudPGtoOO
RIYcnOehN4crHmXNBHYdjlNzL9OapY8MdX/QdXofDyFJsDbyn3Olm8oTSqP/RFEA
lkah1tWGt4Jpwk5nILbGwLaMFyV9AZ4GmkQL4Ia9sw0rcLtgcmEc/cuDLxVv+4Tk
GXNy6wW2gg1J1ulmo/I/4suuyU/XmR5FQgLVLAQ8P1DGePeHEx9BZGVWYnv4sAom
QxHb3FSxwCCfSHXZXm/b+0Nrz3D6cimgW8atf6wGYUH7IGUOmr99OqD8CLJ6ESZg
h7wq1rO1msg0zIBk7qhw/14BZGHiolLeZoQDPKfFpm8/5+jWIS9/ZEZuiHkyovc0
W118CiE7x5xts3ydt27/guUhbbdHPL42fuNVI9wN3Pi35XLiKE+jT+0YessYdatE
ZtTxpdxTyYOmiN+59jX0kgxTsdWMOAyldIOJd+dR+KEXwW9lV4M8jqaclyC1onUW
4pZXByof5kDALOfTCXz5WJyuO3luK7jZs4PyM1EqwREb5/nXu370Pc3csYaTI8r9
t5ShIPHSoPdqywTQta121jGoZMgnHbefdWp8PTuBMIzfDuKMWYr3DEBetEgicV17
K3pFJZSfvzT+CeER6tPI9MtgwZGUJEr6OG2R80eVNO1kac3B56SJznek+DgNH/wn
k15E6GFiYp8a9dZ+ZPfmuYY83nG8732RlQz0gwE+E5mfcv+xGG3GBYsGRV5hJUA5
92glHEr1RXVU84tWi0Bu+lv3r6JtbpnoOyulnV/jIUf7y+RWg61Zgwbbzs5guKBY
usVKW9UYy5HKfnHyPRImsxcEoT26y0rB6Gnxb93h5hs+RwJGRpmnb5i+K/INQBBt
CzyZ/D6wxZwUILVjtsOHuCDX60jA+QCfCqY0n9Zc6d3O2JbYviVwkGk3H1I2I2ia
CxwZ07aX2xycnxlVDbW8Ncs7IJ/uLEdiQGH7uM3S3jK3pF+op2fPcDGuXjfxREZE
a7EVRF/dPsZpsAKW7O2GMNOcrILtNfZ9IK9jtO+C04pFkCToFuCZfbbDiuDPAZ3o
qA973q0enTa3tvMR3T4FnJhGe99FpdDOehJX09CyZ8NLoiSxEaw95O1kjZiz08L1
bzYtcU2htJMLN2xTVRvsGCEn4tcMKFHJOlmFwGCBHx96LEbrLmpaYkeWRmO9Nrij
oPE3Q6X2I4dtJqihddhUESfa9j9UMLLLDI6YRhPf/gmfmbWysVWnNxq4ah73GPBm
u3IqViY0qNOH4bU+r5yjj0h0dk8w3EqORyyKWkXL9o8hCPaRe/6jtXUD/pmSHn1X
qH7A9aPWalqOG+Wr+z4GnFFzXA9LTzKpTy9Ns/9RwX/k6WjhcKMApcKQ6bk7tqbG
l43PA6Sw90mPeoFnT1aXwLjpEhhG3X8ap4EC8bh6GR8r3x9QnuBp23vhqSI0CHT9
DJeYY3sGfExdzc1DtXSd7/2z1R6B2heAui6z+6ukLR5TwW7zFCHdLisp2vvMvgyx
SU8P2e2N+f7jYW3dQX5DnqEoHUQMaVoBKoR2cYbEjfUSG3SVSjyxZluXKFJveHoz
6bldkTxUtMl0eCsfsRRpzN7JgtnizJVF037wri912VbK4n7KwCQkmwAdqS2qlRVo
e1VooG/6uliZnenQbwGmMsE77IdXkCmghAuQ0nl/qkG4vQKgBiUtygvYQZSvapAI
cckx28iDDrAASeGDgA+5fkwB1jGkuztWyg5GzT1Tdaww6PTKJ9qohVPONQwv5+G4
chtZdOeAJnynRnYpLgo6M+Vu7V9+JXLCk0f9ZP/HI0Qr3Q8pqeMNVu3SH5UBZkcb
PMlNksugDq2UPzRUa7nSaTw/6xoL0ZHw28XazNIEcFvdfcAhU69jYxiKeg1JA0fS
yMbkrSl0UWY5aFZOgs/9RduWoW+9qtMGrCqEl1oWxgoSLPQ3n0CL+nW9wbj3JvEb
nWH0wujd7I0FlfozActO9IC9DxTkMBvW9ktXq1cWI+/RI6NaSUSgqh9DrQrqT46b
d6Ols8mdfg6vbEvr8N2fM0vKIb9/29Iu2/3uIDnvUCM/YHcMkxV8uM/TbZnKEICS
tYMz+YtZm5WSJFD6zlvnFYBw/DfjbfHddOKKeYFrvww2CjXy3rO2Z8mMt1br6Uty
ZD+ROH9FEAg69deggwzzxKjg2FeA5ZQXhppCDMHsOqg8D76C70l6frXTbKT4UmVp
+bbOI4zMfrt/rWdD7C/wQQT1S4Sb0QfVm5N0AGc+iR1zMn5Zlk9WO/jlF0aS1bC6
MBPJmvQhNCyP2+SFdKsaCy8UJmSM5k1Gwk4UPlIDcWnXms9zsmo3DVxqlv/iobNB
zxhdEkpeDQi0GzTqy5Kg+2Lem94FhpVEWrpXeKae41fUKsQ+IA7qaF1QlsS50d22
0ITDvIu6Fppi+AV5SBJheKCJmOJHZTp9l2EP8y2oO0XhdGY9X81XcT5p+YXIEU4r
Z794rhjxs+qq+nZG/wqB58eXEGd700r3UnWymrFxGh/IjPGgaWXs/vLrJtMzyCZW
5War4WSQlth+EYAy8Xg7h1qy+ak+wdSvDdfX6r8ATpoEZwjWPHF/QHzeUTwSYjgW
UWAAHXV4tvCVqhEdONaTb2GvWwiK7AMql5Pm9a4V1+Mg80enbTfKskNvl1Q8LHMd
je9GgXJIjQaL3qdngxsnrG5a2gc8mGrSmisuh1QOaaELTYZm9qiue13qxoe6FI5J
3pYDxJ50IaScdQs+2a2mHvynQKuRRNAYtKLxw/pfCfOox6kA3Hq98kXov3OtpXkG
wPEQRAxwE/FUcrwYoKAuT8pKnQr3lYcHBNsN/JlMdUENCj8tNOuFOslLR/tMXHYj
qBuLDC964sks9BsQur5M9sVK4zJT+GdfCupk8E6cYNG0UqCGaDQNASwHqQVZC2bT
xpKOf1QF06isVNr8Pu+A8kcrNl9+C3Nz/xiiRX5X7TLzc99mFoYaNoC5Ibrfdych
thLqp1wTKmlaoHTgT4wyOMIxOTuiXPO8zkMAqsRbtHXjMtk+Ghkmbw+sv2WRHwbf
XHENvr9SNgpjocglbQevBWzTk8bDfYrTAUrnL5cgXWoY5XyGFJL/iIaQevXDF3QJ
aqZ4uSU9YF3COGEsq+wr+hb2MOnoiw6g5fAyGSPMoMATDe/AZQaO1fJLvU9gtpkU
6KITXGYmr213g60Tgr1hU93UyQdoiW9gFh5V7Noxj3rIJ+CHFcxDlep1pMHlYSwC
7lY1kEgGhlIUWdQcFv2VcxzqRLa58YdHfKjXowgVH/jTwyQiytGMiWf7NrqgZ+0Z
6i0QcI/zMsBbKP9lrZKfYH8Ryo6KXeDnN8Aj1eeG4GCJb1QswL/y03Z1MbToLnSO
AKBw3XGQvfTodabOq8tcxhLgcGR94lTIamttsag8a4FN6TDnPLcKAvhhnD1p0C3c
r+d6IszrTOSq8ylHj3P/kiSI7Ct5kxtsVl/q/xQrl/fUR2creH8G0nUZciOeh9c8
e0fhDpuTuKRuxQmGYuftI2zvpFfvg+f4LRKh1K1RmljXbJaeXIb192Tf9B/+T1Iw
txn0R33b41pQ1OraB5QCp44jeyYSCAieuzEM8sDmDD+l6ZwixGpUb99pXDZkYuit
pxgWmLqjFNNFTzvMOr6D+ve+eaHjerqE8XM3eEcf941jAhhuGVAWCZEclFVU85Po
ruy2T+Sf7437N4QHosZyG2X+0VOnCivE7O0fkZl7wGc7pdqGgqlf7qVobypB+r20
BrEWm6GZlmPIvxlnITHYSF0lAgerXHFhnUiiGz4gtD00cJoFl2v/KuKX070HLu/R
1B9VdSiqa3DdY4M6vPDFhirCVLaGLs7ZKhkFva1RYDFWeA0L+aFL9fOQatnuwMFD
AXcJaqoE0j9Z0IiX8IqyAMGmP6ZYtm4vfur8f7PfxAcVNXn2C04ebhzRLAOMuNyd
/mFpCYqei/i9g+oWxt/50bY+7WkhzdbSKeDAtCtbR13xW5HXKBlC69sT1HORqc62
6FbZ9AX2p2cARoeBg028sJfkk/MU+aeRDS6GtvX73BDkFxf96mgnqkG9IVTHiGd7
sdxshoNOUGBtA7xQzI8oKvjin8baa2lDqfzUyKWoxbS3RJo6vAehk/KeC3T9JPyv
/AVng5pOqN3SsnUZN95YuRpkrCHWkLHnrUTJhz38Jj70x/Fc0XRGTcyDY+FNvqfl
FOLMP6lirWTmoQU/fdiP0sDoFr02e+o+EA7yrNaSsrISOiwD6Jx6NxxzQfmwYrvL
RZeiInrrbzAAk1+CSdm9jLCQwyiRVHv5nwKJjGftnSvAvTU4WZc8tt7q+qMrdNiw
iD6Q5ZLA3ABA7kmh5Kky5T7RoQM19dJ0X8YIFAe1o6yZ4DjTNP8Zq851KTirM9e0
xLJQmzumfkNcwtAWvtD+CecdKQAyjDTKK6U5lVFWFwh7E6pOiLCIRtDyjY+BjEAl
KNMjf8GoX17OVKyxH8DJnCVzsN5Ze2pmGgFl9yixrV4J+4guIgZ5T5fVBWicCw4T
Q4pb1DXManuh5Qpo/dJkAZvfZPuosKyNEEzcqZ8L9NG0/zlnq7i7LNZlrn7+siXT
S7xYmSvHe7xMWxlaC52dZc16rN2CM4jScWDBR+rNhmaFzxagE4CAMKFAtq9EdOAp
swbbcJvpp6eBK3Bub0kckF2ODBiq1txOIPJ5Syn8AViAN9758QVM+oApr7mplfVW
mfV9qtGRvTVilNLJqULJA+t/NvgnATUzNMAbYoj9hs3dWZdL4pdQF3IAGt00aD6M
1K7jo3U29CwTHEvm18ZlVEwGu3A7mzzsoJsJOEoHhZhjmVRW+jSIrJpTArPyAzkL
WIqAvPO3UMoetpHXGP3y9DU5pQXdaIVL05Bn9Jw0/kepQ/SNaSpY+UVvIrdmO56T
f9okDs/DQneieldTwouzyal+tArdXAfpl1fi1TyNlAnV1XpJurjzwSaQYgLM6nq6
G7VhwN/hDP9jNC80+ALOody05PZC9MAzp2H4ULvmpB+K5xP+78VBE47dvxdj94mZ
g46PsJXoR6JPbBbVNnbMxfu/CHQvOQAdUw9m3fFdzIb47/gf8YTOgpozyo2Id6ld
52lqX6S7Z/Bt0Dkm7ETlLvhQk9As6xU7UNaYUaMF9mBzMipNjpkIDxcm4tasRwoZ
iZHR/j3j536lZA73ZnXu0K8VhFb8aASuXV8w7DB+ez6enpLq1k3yZG6f5ayZH6VG
4uwX4roOWogQuCOvXejkNsX9xtFRJQPX3PWOQyni14h8tvSpKfP59ise/duJPcpl
/goamiK2D3yL8DVXI/AFq2TESOogr8b1RkUfP1k56wKXgDflDgccLjO9xihoMLAS
QzI6swvfIEZlpxpZazoNdvsZZ1hG3tQw1kk4XDxdxPoh5ajQvS26AU898jbyXJ6y
hX6kg5C9RvACrYp3cf7CMzknSYSf67kis7yiIvvRlGRSuNIxDL0oLGDlY1Y3/r1V
LF2VweWUbWTcdAchBFQ0zqnDITLVppt9XDcoPvegrgQxax6AIAMV9Oibl416FeCG
ueE5HaV/skdJB3rHx6EKBZvgM3CLDuV5tYWhtyLVp2zjTl2f5AQnt1eZhmp/Xb6S
Y8H9GcB868OYocoPst1BrZxi/3q1QOtH7GXLzjV1P++XOoGViLRBgii4KoANtZbP
+oc8JcFpHqLrUEryBKVIMbQInMzpdFE4SnMCN+2Dj0LSv1Tfj4YFrShnKyGZbyWe
/Nzs7h2DRqU4/BT9vKdvXVl9LrQoqkBnblrUcA2u4prR/P5DE+UBRowqEpQTlPx/
DhAGd+By/ljpNtyKpt3k/nR5D9dah7TaIklZ8gS2snGzHBgI/0rFwbDJ1cw3naQe
kiX2YM/HJCA2LyCO7/gZqE5Cms3af3H4SOFvyQ9icL9YvKf9yjzEPztmHnbrBrwr
6qm01wyQHRPyEv2jXFITM2XjzqzGw6Bg/f62cyIw143J7nKrxel8NmeVtOemlIAo
pJg9S7bWb5t0527Plt/k1iWMnsX4v8aK2iyyFXleRSIA6iZS7np1yh+fa5HhEUvt
0x4STbicSY1lMc9rEJ7E+rGUz83FMJvVsjDwQfbbCaLxBD71awGdj7kj1fstUQgn
CyKtgbkuGlKsoVGGrdmG3p3pKkC8Guf4OZAjP08gWP929bDgRExmoBAl7JjeL+Hd
ZcTVryTUrjhSlp2FRejGIWlKmWDLNbUkAMZh+6WeczNzHhFUnxeGR8rV+Dr74FsA
8nnIcOEJ9TXmmYix8G5Wpx2xH6XWKinWaIOVpBTR1H7/lrwjhJqTGrQtZasV580B
cL9wKE2fS0xUty4xMVrh+7FDREl0p8LGGc57G7bnz/44u14DpRshkz4Y5kOgPl/N
2wGgzA/OCkzrg1eArkRtcsLYwJpj4W7+McDSlulgCa1ty8M/zD6Er64rM4hovSrT
Sgn5FSSpVOLNn2ouRtnWNwDofvZ1wwReSYqyMU1CrNMe57vjuB0qcR5q0j9ghK50
Eer38R+52XOH9iEN8P8M9bnKl/Hg+sp4jgOSjaW0RDeTUJMtW33yUQEM5tkgTEu2
nEQLt2H0meKfZECpKFv4OikgXk4WHY6lPLmTNbLlE8Qx7pzaP+7EdDgtY64egBnY
mGlssaTLdfSBUhY80J2V/pg8pgjjKMQZ69NNTp5HxUrmLWkApdRyWahd38b7ASOu
umzvwkV6aTi73rjLiELYagto4N7b8NAsMFfrkGl54HLOY9Jk7TaorQZWJph3U2Ee
aYrFHs2DY+jf2w9g8E2ptf3yq3EGI48ATl9NsAo5u2IT9BAHpA7awONHtrUL9hex
Us9YORFk9sYkBK63UMZ+oKOLQdor+WEVCYWEZCnhlYNHEbJToifNVhKY+wXUJXuD
60dqLXbrgTWpiAaD79gcGNnKjYGbEr+D/bkoxJchupthu9+wpXqqgLR5qKmtGtNw
9p2ycKverllnE6mhuSu7LBhR/AXnHCYDw8tCOziVRzmHsUFDJTAAOoufQhjQQQWQ
+CBVhAqIj1VS8hKOG620xUAS3mH/LzvYeJpA8l9LlifBC9Hc2EmWo49LhOlAgPA3
94VQN1vMxNq0qNBp6anVw3RHq1qKjnKzjSlezXBDbi6ORJNyvsn2oNX3+DOm9DmN
3XVNzg4lI8atlmqbRQrlWJzEAF5fAgAn/TQ2hJ9mKwa/4ctvBK0SXPpm6yrj6YFw
yXO3f/qRHOcerQNzjiUy+yzZM0Edblk3OdzPQ5U7S5+jX4sGmUIjf2U7sBP8+ZtB
7BrXMC6kz/IX2bgPat1nBW0P0K7Om41rqoUQF9z7qkpwb6M+YXefWoCExMbb+Sbk
IVr7sc1P0yXcBtO1j8GMfDJT2tLYEd6pDXeZM+5rXmUfBqNOHOMqupvkMwGtkGcR
0ETl1DwS7kwOMZQ4MhSG10bQgHnTC0rxn2ptxKWsuEC+Sfnb8yT16Y5x177V9HWs
cbpqZcK2S3FAILm20BO5eVW3p8KuInSbdtJApQrBgbtRLkP0hrOyu8hBZ/1LY3ie
DnUZCM1CEHFDHaIZYT+VbZ4RW0t4EXHpvLH/gT4xQTVJ26lX+IjBbEJ9yEOo+HYh
PujESFwsp9um9CbL6rAcAKOQXgJ7rm5/OC4KZ9ugpQ3Qne0ozQ5XV29UKiHJzzWT
s+AqQtcB3ecTSLJ8jfwycZraUv1XQ/gdGc0mP37Pu0w00lz7CBzJE+dZDEAe/ggh
Vy2yjLeuUQ407eAjU1schJGUi2h0aUgGgBlDmtnGV97Hfh54qEA+HLYX/Xe/SW1z
k8zcMxrll4GctP6qaJAd5HIhLuhikFK4pZC5qH0goVjyO2sMQmMF9GopqLI/9Nsq
C6atINogwJrfFr+r8PjqJHxvefCOuo1GIkuO8Y3y4PZv7hhjd1URUMxiU56LmBm5
IaiECfEoXCYghK1+Usd/bHcSHAZmzq6/89hURbb2DZbDKigZ4mrsyDnSboxzqsvm
2nQZ2DomnaquYUhk9flrUpVTjekFNtpYSBxiS8M3LbJZPPCd8qRNKKD9DG4b1y8j
nSDapRzQI7C8T5JM5er4VbyX5B6/LCXT/d0h7lnGoMwkXb8msP972T2aFCRossrV
FQWcOcE7JpcCSE+mW6mdrxvfEN+iqo2Hd0I7j9uac1+jEf59xLvN08D/xiJZHMYT
oPcbbVZq8UHC4Lmt/n1kDfsHiwP3StUN0SwWxIb+9SU9OTAhGXVQ63t1QzbLzaXq
hSWEbMuFtkiSq8CUOKqovNZIaG7H9ZuyJu69HQR19xJnFG5Odti5i54IJQBmq1pW
xRj41uibCT+uBGl71GTuIq+m0dsbkWwKCW0MJS12ySG4SAqnvc3UcWpE24agXRjm
YVtfgfEygHh8r18lXYuyVniYi9fX15D9ORYhl8d4IW36n79JRuYn2d6afuus27AU
+8upAVJARz9KTiZORZFQs/3pCP74PrqdxGbcKGwBxZpKkYv7j2bW0sdWCpFvxtXs
UQoJ0l+bW0XiDw/pLwkaci0Qy7ysZuRyw9LTf5qbOaol/6GQGW7XPwbVfXi2PdzQ
31Gp9SjutFy8Iy9ahGXSLkmlqiBq1qOsR7hgof6aJP3y84dQgndp+q0YuSFLGn/7
pxDuk795NB6TL6y/UAB5I7y1+zF8uYJ4AIf2gpcEfo+1NPgwgUVdgeHO7YzbGVIP
zGpeIiCbImg5lIHNeBygq9g/VTMEsS9xLp9eLe+Wis/sHq0GuX1+lybV5UxcWwZJ
a7r2KfKMx+iTh4VmCMggCqKbfNHdorsi0plY6VjzZteBPPst01/NvkhPx9aLuW17
U472gyzy5f3nocL4TsOH4jbDQ50WC99G4MW1zJaSb0B3dilpYoVH1y30BDhTLsPx
J6RiuJ8KMt+v64aJPMvghGgU/O3nDbc7bhbx45xwJeTGbb4QdKmSbLDvlpbOfwZp
HReT3zmit6pVGUaFuidLuEgxyPzQBn7pt3IVuAkUdDRgEADv2poXEpCosjGyEjem
QPpMfhiW5fPCnxDQCpITxIeXt06jimqE8FLQxdd2Wv/cpa7hdtUQvGQ17US4QVZ4
ciy8sHiFBUyCHgdcRybJeFUutr6LXcUMbayYm46agt2iklSsdmU+cyOkexRWVf0f
mKe+RzoZuSNTczVbCNqzKf/z/THyLGhsWa3w5FI8QSEFfMlT6a/t0eXIfnJJsEor
5QsHyXhvhjoC+grCnBKz/Rc7/6IL7jfyLrmvBa1/ilZ8szGKaWD3YLqj1DP8pwZe
iGrPNwupbJojwh3LPd1DgJUuClr4mUGFkFCl8whHOokD65NM/e6sB/y7PWHe3tgQ
hFZC4ydChnx0S5fJEO5gQJjpa4cJbNi+8s0ePRYPxZBNY/gGeT6ucACvJRv7147e
xM8xkfvuD+GEoTdKHTo1BNNa1vP8nGnoeJf5y/gpp0JZJ++PB9WQ2j4KZ5PavvGX
rrnJ5cqQBGL+QCjfIV1unXHHHA8h4CNOFDbyeG5RrhcBPf/geIR+eJ88ALuCIKVM
evt3INOt8Jt87AXL1W/kdRonNlsc4v/5MN42P/3MnHhANwz8FwZurYbKpqk/bCVD
pyRG+33hJZgEzFnlLp21A1P6dp+BOWHaPGy3rkJ+EnGtPDdDHepO2+99WruL3M+h
r9mA+RlmZNLlG6eOm3LzZs8LCxewiRMOhtR9z3glo6CXh6h0mdeInbXrXnBk56Yn
k2wLT8YAu7z1BNaCtueH9H3i/OilnQCmN5HJ1sS9IVvCc8WLtGk+pbo1H6DhP96j
guM1pmDXMwbOzRCh6ZFxqekbTFLUgGHeA86/yh6diayvQ8mCMgvAnJv4PRAEz8en
xElkcYM5Q2FYGrglDHP+XMULo5rJWFJPH8d7A0+8ZAipdtH16sBl8/RTNYznELun
Y1uU1+2ogHVKqwBBhdSRfHw6PRpqUROVrxejzrjkbZjk9tl/28bHOArleGYPR/1Y
IJHBZAFYtIKwNK6SsGgDyhnYwPqJ1av4x4wniKjjvyzTAvtorrNAjfohQw96fgp9
vf0rDj7v6pCAmRpApTT5ijPbYeRSRHPpHs0ecObMXqqwJ98atM5Pz9DhmVoRhk2h
v+SBqwNalokmFxLCo6w/7ggV4srNYZRPad31/LrvqNplS7lUsuFsOcJfbwsCsU1b
ErIlHWUQz4tPt2Hn3tLVSNsA6NN2VCui5K17lNv2psrNtnsUxvIFLGGP0xeyxbFN
pErZLhjXt4b8cT5M2O5RIZQ6FAy+65l7KTjx7aqtVr2ImiUjs9uCGyrWNB8jhvtN
2aXe9okjiN1x5WQXSTWLNVq8fVjs+eN76OrpOSKrC1C60Vp2KZxCNaYptfQq/slB
RC32gfyc8PEt2L2T4dcsXwfHTQe5WtTk+vHqjHJB43YNHC3nR/EXxs5JC16SIjgy
VAtrmFkrUEDzBO1RQVPp8wMe9GxIS3lz9OHI8JWo++Fr/ddf4+hftsgbcl2AboZC
fieFXXlSStbrQr+NupZ4EzoDTfWdw/PFScSwHtcfcy+pSzIf4SzeI52VFN/j4xKg
UTKyTL5rLZwpsrWKBny1Zs0+NpCLxPEogREDvlgUKvdblfzP8wBv3C8GEc9MKWwK
sptFhHB9zDSRgvj8yceTtWiyk/6rQ++BQxgopw/K1G3GTgWp0RGp8CAYBKWvPC2H
HbVKjOdCAC86+l6O1PA9gtlLDqykrWk7rYN+l9POsqWXhhIRtsNQ/PBzOskNtN19
2rlEIdmupA9YBHJqBJV9Y3OGziL85oWsnqVtCdpBmr12EoyOP/Kxjww8cCmaut3R
RV0+pZbkI5WaWodmCFveA8ujg9G6yQniVHZ7HnKc2WJt8+WCg4cRLS/HGyApIxlB
PRWaRBQZdKnydt8YtPsHgeSCGj2xufx6iucqMmscXGdvE7VMbazw240bdqsRehlU
khm03xrQUL+E/nkN6NexA9Xcp0ZtIsfzQfBzsh9rrhHqqVzxdkV44iAuj+2FIgck
fGt41yjK3TZIFaq4rALWV0dI1rUiiBODPs7dvc6dWQVfFmWV9mUyKGkIu3aAWtap
wxVH7x6mDvss0xDp92ppHGqHodPiIPj0/ivBvmBqjplDkFGsvFbV/lFG+f1lQ4VN
9o+vVNiYYAK0JBtbewsxjCOqTqJFByrh+KG9TcoeSlvCrb8zwpGufX8K9+2PV3Mx
GDruZnQ2IQQev0VlERFRCx6t3k2rBgGg9TqVedcdFgr3+jZNWghTajOYhbMdbap1
7iP+rs0Bc1WBrs6r5TmyG1Ipih6oUXCfD3Kl32VinojXdJkct7ofXBcWte39N55n
cJtOjyQsi17l/vGddHxAAOSTUyuqdUzpMQAZwKdZzv7QLB5gfyGVvYUoDgKh7SV9
TSCNIkzz0YmoQcYF/R5eMP5aQ+9Xhb47EuxjLKzNa1d+Xmi5vJDqlBQ2exxBM30E
aMXt+z9EIUzUjdrw9yaRFzfaEDaTBp+nqhv9FbSYFe+SY7m1HaDtwGCklywFpiWk
dyEehiRuPwio+F1cKwz3ROXKYBd4d6fsyQYjf2ivWrAIIhRcHxaNaL3u8kqZCsgN
2vQYj69Qm7qvysosR6TXH7Kdu78rHoFsLATvQ8f0WKDGMkGBAtv+yJgTDkSSvphq
wjYC26nXo4XC+lVms/M1WcdzcR3KLgYHdgsk9ZGjX6CXdi+c3gKoLIQ9t6G0aqbn
b8AxzQW1e77Xjw24PAzObPH+N8na8iOVfw+YW7ovTuxt0plGD/EM4LZIfj239/W5
ILSjEZqY4hZRVx8nJWq0q3KV2g0J5N2mhbtfDnpTKQOZC3IA4YGnjKjaI6yM1V5D
OOU7Vg2/uU9WR1PXUVGj4CrEbgniA2zqE13AgRDzaMpXELzWYcb1gCKzbSbSIzqO
fBIU0+kseqJzdImfoHy5x6B7inq9Gos1Dl+LU+Ej+oBJeB8OVwg1KSFzrq9twbMm
0HtkY9Do7kCrLv0Dn7QQ5IoglxK8AeTkSUm8ocMKLS5BdceapDqwIHJQyFk4M836
Ff2lKIETSssYP7Xesw09OQqPLqFIPImAv7ty/4WBPqpcwk/PW0HxmasEONIpwwrj
4Ni4ZpzlyTR0iQx0MFkbqguUdgcU9y1SCzZIL3jBMtTVTsnQQe12r7sO56XPctpM
DaRE2XjeL2KmDpPapT1aG7rEQA4zQGWp3qbKLCvv6+yocm5ujSYBpNyb3ZUQ/2ZL
Dzwj4oNf1vp1FyVz2g1qc7F3SoXcoFb9KXC01mY5jS5NLL33DyjShrsdB/klC9kK
SZu82FBTdjffkJ6fgKnnqQzkVT75z/xSaNY4XHTvrlTT2lILb6npbA4oReZdVT13
vRUtk6PfsBJnk6yzUDDWupVUCQeC4idaT/L7xcWkmqTtYuPZ6y/G8dmCBRrLfIN6
4RpJc42XX23bDDdt6jPw8+qQ1nw16Gkp6un67ezOmUBbelcUh9R1fl7m9srQkctv
tSKQsXOMR9xlHo+R/9ha1rhHHUmnBtKubn75PeZiFJU/IHwPy9fqoW8RjqvwP4cQ
iqWp7IKwJ4AZ+Z1GFm8npF5iNzwOIhXSjP8qC+pDeFAo3P+du2S1dwd/uF/1uX7B
xPSglgnkW1vy8daZd9dmVuO63PNrTFGZuiXlcwRYXmTNmr8Spl3lawdn/3iNm+Ca
dodmV3VLs1F+yuJpq8K6E//ikT8BaOAdPC7EVxsPoDVC3fQY1nq45Zt5YQ+bkPW9
WZHthV8hqEQK5Pkga7Q8g2KJLkE4h0jjtLgp1ycmGD7FtZeYEZciH4dv/GqqZ7s4
I/pp5+BcwWbFfQa7UthLmwwfyuElrPb+794mhTe3v8G8Kvl0dfPlr1ihmx/RUY5T
q9YcluXuSQ0NAxj9gMiUwxO8bu8AHlHtaAMMq5KxipHmQn4zkjQV4gLNqKGHGs0w
zbtMA2sEJFvN174YODNtMcVBrzzE2HpqVY04nzzygRXPKYsIGLUYnXFCWhnutKxG
3J4lcZimgyHs8FCefqb+Ke93iFFR2BwobtMcZKX531Pc8LRZABe6bToecZD+6BFI
uYJwi58wwM5TVDL8OAItBDXGUFFqxyz8s8k8/qlQqVes3BahvVhNMFZxMsIqo4og
j7Kzi7iGvfjt5mkrhsJDHaexbgWNyfy2Do2rpXGRneOFWWLPOAnyzjO7BiqULoKI
QkkpuzlQNvWgCF+piEq1i6QteHnH6CAmMvcZuOu3yOf5eK8EOiJseOW0InPLJbvq
lCbw23YuUKOURkMr/BG43IcPd/WBqJwfOelGpGuxKZoQzBXDVzNuTNS0u5nPVrfC
RwU0Q5yrf7FF2cxnSWktzLlkAM6yqqI6YWlVaiHBUb1xVZXeP91Q3FkaKSnODLME
I5bwhiTkYRBCL9L+ugwhno5E6AI0c+K1f3XyoEXHclQibWsFTWQjfP1eUZsTgkkD
bTjMDHP2OYKe9jhVbzv8LialYE/3NsrEbqehyKv/773vSi3h7/6av+0ZA+qjHyAb
WxwgtKWmnUAXewfukJo2ZRJ9SYK3jntgLyQYnoBgomB581PnrfAFhk6/kmmrKQzF
yteAaQJiD9Mqi1ZQRfa0vpYYkMI4kCku4hFYD9ATlE3cKpcbqxA8nttenqWDhc0/
Eur0E4EJSgmZ0iRXjTp38Q85NZNodCCbrZQiK/gUGv8e31m2isiFdKPJwcxygilf
WewGJ+ZdBWqS6AmZqCNDDoz8GCGAKK0hG7w/QuKuVa3j3GFVwKG95y8XsdYD2kZN
QaDGnzpU7jErvOcPDqdqja8aYaUZMEkOxjk7xX860nS2QNsAw+nMfuajgzWBi43x
J04ThGtgH30jlgeqkJn+NqP0kkwwr/gjoKLoCPFBbZb8GjCGFumkGRvzwQ71S7aM
hbFUP9+9rAL+bS8KTo+VE4zn6/H+gKKbCfvuZxLIm3BwXPj2A5zSyhis+9X5Azco
MZvOy4yop1MXjlAaDXYHVNP99uEm1g4Q8XEvK/TvGyOyPIyJjp8vXS+tmncHKlYJ
GY8Yv7rsWFAyXStOt42mTG+k1Mlo4QhUpxvJJlmbl93M4sGOz0lLHnH1dHzAMrNt
Z+50O8alOr4tkLOaQT/kkw0iVdquoCyeUBhJ+ZfcHZZb79FT3SwQTkoQ/bjTmZtT
qLKV14BE+4U12/RbIdp7ubujtbCMO1QI8FdC+0lr6j1NFVN3uARQmofB7JVuiwdF
4uiRb2qmEjXGhfh7pG3HBVidNNX0ko+NciUCei/tHxSYAWegggU8L1rgZInDXAoe
w4r140RJYxJgcbboSpMEy3PN19lTY2Y6urZVU3NDVVmz322Nf1/EbW9g+26Cbzij
mh0Kcx0QNtn3U0/KSxg7jxivCGEiGOFQR9F5jNAYCy1+d0ai5xuTX3SUa6bCtxq6
G+RK8g4wzj6UfhDEy+CS6CcKdUhxNO3/CJSYObi3jihV/+X2ay4N446CifPcpdaP
NJvcKZbBnKUGdvKIGRHkLN1Klici83ICw8yE/u7riQfsGRNCS9fz5xKPbnI/LsWF
lUSIzDHYcXpIwLVg7LNUyYON1r+68l7BWw4TspGXI34NNwL/IjyWs6L6ZnFWYLpP
9G0YY8bNII7XgTTnMENaRV5Ph9tJ/6hxfvaD93J3c3S9d+NWRGDACNCtHgebKjF9
KmDz7sysULFn5bWNSX0rI0JEMnmPoAZSMsklugu43FDF/mXxwv9RJoaXX/qMuJll
tby3XN1khrDMnPaIRb/KZdg6AA7PVCIJdWIRmEVawsAGS6HijaE71h4FAsDSoPEi
SNzyacijkxONRmqfi1Dq7+BcmiArLCBQ1j6/Nw2bLNfMr75moLaPrhWiEWGG854I
NNX8pxkhL/Q2k/c4pxNmxp4ayUYXNLVrQGjhbBbjg0FkcXtFZDq6y8h2dJmDsvRh
r+dvR5MPSFF9+YKZ2UESMz18SnFmJFR2btNlP7Z7hcaJTsh8B2ruS5woMYv9Xzes
YlNXmDBI9gO37JwTeb+3djlfTf21tD1SpCPAY0V5qlUHOVGWEVQDOUlR6Hl3q0ld
BaDS/nN+oz0eCnH5IWtbWgg8erpp+yub1y5EkRpBGtdCRP6UWiats/WuPLTpudXR
fnBfVltGnkkp1II4C6O9f56Q1oPCnXjas40qA+ilZ5k4dWdQjslA3yWgDcaIKkT1
hoTuOs2pQiDndUVzHETaYMdQ1ytrn5hsFyr/9Rff1R3oWbEnvfJvseNV4TCTPMie
K2YnI10yS4tvgIIOuArg44KBGVJTVNxKFHKk55YlmtRuAzcIKi/PCX15SORHLyIa
L4Y2IeEIHU8roEbEvZG5RdtMrQ8/NdB9388lWaOCHJ2oo6Z7Pnd9VCp3A9xZStA/
GBM05xY9BgdF5K+aaVvMDiimNi7FPkINRRsAySbXE5TGkyJnRBG66m32awZBKCo5
OJaAJxhPFsjS7lHQyZXIW+/MrNy+aCznPPbn1oVIJcUDAt00FpQJ/wj9VFt69beX
44s/HfseeTdG30QuPznzfKx5NrI0LzLNskG3chYYVA1eS/KualhPhnCpma9rxsNI
IPaTbVLFC4rpOUxkT+TRBR0R8wLppRTNPXwI217UFxpiP4Nt+rumRZV52jXMg5GY
vArC1B/9i2Q/FC/d8ywx9l/J8wdVYsNZUKzk59dfkyN71zdeoVXcJ5VAg+hNoIoL
caVzjWRmJFwSyWhR10ikFDv/twuACwy0+6lT+7gnW+r+csjlMAMZgWxEkOQ53wm8
eCgEyosSZevybHIylg7n2cFeZzrIXPxElgsINPRlvd+gtREVhH99WREdc7uN9/4H
j1lhZqT2R3dyeuPT67SJG/5k+5mBc5G04B/oyFIxueOQGPsEsBuNWUrn+S7j2qHP
ouh9EDkTPH45sz8ihlnwfvUGWrrtNdvw8Ar+96nZmlzkj1F5Uzo1HMmgUXdtp0Ri
nqlqnSzlgguobPzT0Q/EMQjyfkZfAfs91HAqD/QcpzVfWnxGNDwPvAoXwfCwoi0a
3SVlZV0/IMBPkk+yClSf7uD8VrfgzA3lEZst3gyld8aqnUzSrTRFFdnpiONac1Y0
OauiN9bJLxEYU2pBduZETsyzaYmli2MXBPrRBF9xXD0QCRSjeKNfjJfuUyaBdk1h
uAQffPikq/EurnPV7H0pm4/ksHWOxhhaxnP4o3k9ZerpRN0a5iyMiMC0GOfx+tEN
SThJdOzuY0uLL6QFHxwQzDl6BItMMbBzI4Cr7nwbHEXU4D5hCmAxvMSarmF4+N63
mxnwlwfCUGBDdyvLvXpLIxnXd9if87fKI3U09AEw91oYuz1l2MN/fixvWIUP3eKu
B16xWMl5Ed+kGmsMr8J3W5aJrsYcaj8L83htEFsKQGpAwLaKOD5bBY17gTu8Jx7K
XqvW7ei18DjyND9KHVeplT53BCkYlV7xfMNkFT5lMGGbHJqxbKDXWENJbCkhlK8Q
de2Yc+uXFIQaErPYvNG5Qhpdet9vA4L7V3RAvMbNy17AZFp9SY8KEOiy9C+UCHtS
Yyu+b3QwgQl6BVJ4Hh5l5kDTqw6tPs6ogk1xVo5/D++mlmieEcS1Phu3JHeIo3Sg
i6iUO16Zg1fNLX3WgaY2uc5iCuJPYUVcLgRoeUmlqH09+JXwUckjbvO90Tbx1FtZ
rEUwIfIYqzO6Rlacp3pCHw1Kk28qWViBzAeGT6TeN/a1+CbHtoFOv1lYbCIX/GaX
fYsSVDzL/Pkg5bECxc5W8PaSfNbWWQfeFtRCb1hqx17pOvG7RKUubC8gJTiyP266
yoiK8H532vpy9I9jT1gqmCC3vhTeGECVjqJp8u3kYGPjXN5ERNzFqk6LlkCHQwvB
BvptFMk3vA/6sK8VxV36OOrqLqsEna6AYLFVbmkhYoWZYPx9nLvHpRSsam30E6Uh
1KG+7T2wOYpWASsgLnyUm9MKxRCKNKsSfA64UnoD7ujZc7/w/5vuqsENdVjjw26S
6pnF/qBVOgcatk/ahpM/FrvluMhWa9cW9JX7/xTMArY/+kYf0H9lSEDLtus2OoA5
kz6ieyKvK9fx5l2bh2k/AKB3mMZVEvK+q590PKxmCNpWfX6cfoQnBBli+BS8iRV6
8wsFM6e3lfYy/8tb4Kthr0cX4WbDXobRsNUaCi9S4odiaIR6mkod4fpe5aqLZHKw
nGIdchDcIOSsaYKKovKzXDhG4MpXbz3EWIQjbyvSEd0eTob3I8dEN2DBrmioti31
+K8xgv0kPTgZxQ+5P1DjkOXGLcZRyx32NPAou+z/rQZjc1/v9iG+aKp+gGuL1hPq
0EAGkPmv7wTmxUo0Wm+5guC3iSe4egoO1LIG1XqgfNsUPEsF29W7Uy/OT7cQs37x
E2/JOxduQRRX7oxCRWgmBVXDMO0p/W90USx1QUnHvk0WhikHoka/IfXVcO9fIu6e
138hkkGgfWl+LmzQPEXszQGivRwjGTZWkBmS202SChSqHR58TfjtM/Zb7JSWg2AF
kkiFBv9xKvxmYLGHF1uP1/zhvCdk2aUl+LVzxninWcsbNcYrsnQ2lGYrXsw33euf
SXgsGScM3yBDomdkwAxzOB2yOdHUYXHYPlfKLYAeLzJfuv0RonZ9Ztylk2FGx4ge
dXILMYrLudZ1v+3d0OzMz/At0eBiidlx98AJO+2+TepKK069qczbyafaFOToCJrg
gfTWL0VFWKqXAY2RRYzpYphK0bSVCiHsvhFX64JzUQAceCFL3q4XP/G+bi6g6B60
9j+GGo8a8gv2qFJn+MMXGCc74U2yU/vew1RSSE4l016UdHVg/fYBi7GRxN7xyWaM
TLy/zp9kHe2lW0/Mv++7nDjfVUarEMu0CMSP7UzgLWTgK4nZnInLB6fhHTHm/UZQ
RXy18cecrxTKGOZKsZaXx3nirgp4g0DqcAv6q6C/dOmVKXkNzYWrld0WeQve2MFf
mExXqC5qCISsGZNqfjms+luwQZec6KiVvbrfaDTtTINZ77KyX/OrQY6eFyYTs3DZ
Cm6qniJe/muTJ8ojcjRRqA/UDdnl0dE7A5WsAN3IXXb45UIPf459qJSUCZCnRx9l
gdrilzQQrytHQqrS3yp8aIJjjTJL41vf6EgMwboQM7QmSZ3Gxm1du5syNLGaunSi
89mmj4wHcL3HB6p6Q7CCWalHj/dq2WlLZw4uPUWtAJeei6hV03SEyC3PRiNS51dt
WlBdKjCK42pVV1cWYd8hwvNLp7Sfb0LdBbKJOR4Eg7mVvJIvbfPp8ZzGLUURRcOD
3BE72/aLHaqEt1//ClY8CKWpwo24/euL6M2ViYo/eSLdPhZnIbYQ7eFcXelBUNGM
rN5mZRyAT+3PrFCRmozdv6FooTMxvMxlPOZYu6MIt/C5ALZxrd8w7i+iRONjS8su
I1J5FQPdvVbCPkHEQ0j5H2ppefMU2AZJvWlUIOTsKE2KxpCC6L1pPTEsUiDXfKdO
zYa+KkpEQLJ/mBrzOqutxHfFagW8xT4OPM3W0J5kjUHyVCizK3CbstkQ9AR3j6bR
dKQvVkyzn1LD86jgC/g+UdVJDNkiizyVQKAVIw94f25oI6svw1IvL+mBeD7m3rCZ
cB4uUeX+o5LWOHj8ANypBLb4Fmo+YURVr7IlP0U5tVa5cLmSGIgpH7adI/uRl+mK
u699yfrJRPc4QzIxucYNyo1ucld5wUIX808iQfPXN8JrerK9N+VXFKg7o5UTlNM3
eXsSK8V4DcOkq3qHQ7jSHNfK79f1YwAmlzImp4soKPzYiDLTcYMVh9y0fXAyNqHT
Nnf+jlVSSi1g9shPvG4w7zQoXZOD9fGsERMh4kTrsStr4FJxNimBmlBD9xEBbseq
Q1n0xijYrhylEC7x+mlHEl5o5/d7rB3ht6ygytzKdJ1HJPpuHM9V00G2hPRSS6xj
YQ5Syk3YeUilhtTkvgttGdjNFHJ7ZUOtjIvBb/96RL7/WCBTLIZ5c9DcjNQoRiu9
kyT3ES73+8/JR7tqTIsYrT0c/Mdv/OMsbj2w8NGfCdDPbUwkJTYp+UfQdimIei5/
zhJpbJj70aqwvbUrZy28oTbCW8TcXy7e63FJPPq4lXet8M+qu9idi67D9JhAtU+j
LYDD+I5xVrpj1yyJvLxgRj5sBH71bteBZHeOG7VpXHmkyckJGSQenyTzZ66ljmyN
VLRCNYDSvUJ0jq+a6SjkNDPUO+2hqMEUd8Tfv5a+dUeroShble+mTcH5MdcqqfLH
ZBH85dubu/anNx2mwUHQNxgFyittwB2rT+inUSPcaQ7PCTdruRdWa3xkO5rPUU7B
oOK0B8xbT8+aXQRQGsgNGWklQXXaMhYh0VgIy2cy8hTgzX3pF4AktKwNv6xleUOS
D6u33ZuHlglv7kkoz7PbaW3TSvMUt+An9o1A6m0ixbUxp5IFX0INJ/HGyyENwNwL
PryPOu0a4Dmjv5EAlcapA2sKP1hzA9RzUuSeJ74ExEJ7HDfYcttRNHYD59J+SCul
UoRO8zo/c0il5Z6B8cnXJzdyS60j49mL6DCSdP60/4xBLzg1iycIk64atEkN5HZn
Ds7wnfby/6/9Q+uILKTd2SbJ9JaJmxJ8UrGLVaG2UJE0GpWP2acnzLerfS4v2W0H
hmZ7jAWJGHZOnrPUzREmCKnbCRSC9Fk8PdxFuauAghZhIsMu8Upa06S0BMNVUEQ7
86ZxtlYtcEOPQwKyw4/J1sNnRBWcVfRRxll88NEmopmT2Vq0at985CwYbEhgMZMG
8QREGctMSxpH2dWxxOqJnQvXac8q3Dt90b0d2f4Er2wKmT5v0V1wsJX3MsujA+0p
/Wrj3cTzSn99mG3ATplyNaq43aJ4M754zirD4L1a8Z9pIHxdhTQ5Bi0fUM8WHgpI
DyYX6Fd6tOVPmrM2ACZs47dw23RS9i2l9c+GJpnFBjK29yo7nyTvp34DfX4epLU2
KBx4/eNEMuQB/s1rRzkRJZZLUMhtxArM9m/TE/X6fXz1XHpb7cpZiVt4ZGdS5u1o
tVSg9iDWJawIJSTZkEnp9UADVkmIue7vXN0eie0WgaN4yod2KqUycPJ2vEIPI9bs
xdkt3FY65Pgi7dEOezTf6rSMOjwNnpJ+ZNlKEAi3B8g+4/xHSs3IYsUUqEtuHbdj
QX3nOnw5QqsvbFWGZqmz8QRsIx4q0ExXirtDtiZ3okOB1t6t5b8tZCN5Qr9J1Z5w
c/CC0tBMmbaN4co/8s8mMS9dM5Co6P00UEQOtJRW1gn/YEOOUWfqvSVByckeQxVL
HcJWEOOBgqqXSuetNujsDe3cxOEvS8xFe8BVukxVgHSDi9cuZ9rlHjyS2/tiaoQO
M7bffE55DRLlDWONhfjGqd+jkP25f9NO5dyhIe7vhOxq2rPTkyx74BbM99pOwZ5x
MIaGZR6KenXuOdgsCM4ZkOdYBWGe8TKf0nNXVrBfwOApZjA36vMD9j49rOYljw7V
KbcwYLLkrdqqt8ZObg4oXJ/Lf/OEH6mVVjgVe+MO2xtgVO+jEt3SipaC5i4nR++7
qBcTI+/QIeNEuPHv0WTjUp82dsOKK6fuByhwhTPNgk7oycRNs3aFuU/Riv/bT/6Q
OHEzC+DF6hUSKVGpz9PdlyRCeFFviN5baFMmaYKos6aBjSJGx1Ed7vLDSI1slEfB
qh3YsiUlOS4PUYxHIb6wC6FKi/7+SBPhUQq9lcrAGY7a+FpuL9/bD18G1D4BeHVZ
6aeylVxWwjBFR8yr6eFNY3KvX8jAgiNTvWyf6NGxrhLvyq2VejHD6ZsMA+iEEqsF
c0HjFXt3Lkb06D7SM8npNoW01MLRHPyecBwn7PKBiK8zk2R2F0UzQdNv/hnWMjzV
+5atD84K3QFw7L02yzmeV/qiyCidGJtF8jRba17M6YumG6wuQEU/4Ngg0e3TcudI
Pv9Ht5c4MiUFegRuT+zYx2gLQzDqaCncA7yzywlg4ueKOmH8tQzyIyqRrMNKC892
t/w/6eK6eAvh0FBl5Bd9js/cF5p6s1REzUJrPNn0saWffDQDPGbRAkY6vtIQL327
MuGA7ATMacJeHKdrKv3eEnIRK26cHbJRpZrCyDhp/9cKyBsiroUpuIoCzybSYsQM
MyBnwZ7+LMECz8lwv+VbOCiwccxgRH4EnZ0Kh7OeAa8a0+C9WM52NKnMXuF5pArL
teX2a8Smz0ool6zwZgbGyGvrtX3SnMbmmgOfNXzW6Qn09EMRTJ0dmlUyIhf7dtzc
qpRkGbHzMycXf00WGX3LQLPDZQhZ2Vefit/3ub5pLqXaz7h8tB1TqocykZmV055R
e9BqvzZJZ/rzZF4Z3EKgxhmVc1a5yp+D+SofY1dpSpwNdLbeUpVag/crzlJaxjrM
qQEOH+bXPNAYtI2TTBkCCSF+oh+8Dl7UBnLvFStlpaCO0czTSS7RDotXXlikfQ56
EJE0Xgfh5+PvV9twbCBmS8GMZbXaLQ1oUuiKvJMxA/lXZ9xHanqm04OheQlzhJoa
zdVfvODoTdwh15BVjiT/VpMI7zrPylOLGyc1UAP+rl+uA84kZb4qMI8KecTsrU93
W3s71l8UbqVnPnr4AQuQJhQZTborA+ucH8lydsO2q02bKV4mBJpKhD2fazVnbPob
OpYDwbNupp21Vwlzdm+3PeEJvLznS/TL+oa5p36CuJ2+M7InNzwhI8+6h0vqDCYM
XQgoxzRyHs9zRlWXLPCz3/LSqWmmEVfS12Uy9tQjbjMQy74aCWWACChcEgWd2aFg
wK6SOj6C1IuPnqI0TUKFsQnhI62zyTNDM3aXg+7REqGV/6rkSTQGSeD79a4R+SX1
Ae9SFv0j+YJnwVlvYJPr8PRQiW0ZB4fwaja8e0tB7I60XLu3EYPhM97DkiWpIsc2
+bhQeU8xgrlkGf5HhV6tR+OBxJowKjggJdZK2+mpP5xJ6PZLRa9taoNaIFY3Rbak
MtyO/D3DgNXkqAREpDq7Khg1lYDihy6XzSIf8ESey53U8qk/eqBNs4pyuNisy2L/
blGj6bDB1hJu+x7ihpi8xxMSMU9BIDghfXkZqHgo5udzN28ku5tFmlWI8JboFVdo
fyOWtmhVpresbt4T7navObPcbSZWcO/E6138MW7ZUeP4WSUQV3op1m4INGi+03YM
7dl7iuTN94aQrUhL7Bm4PSLNZ4ftyFX1ogyyJyLRJuZJFqYHhbx4cjgHhX+13J0E
NtvO5QWD9mEXE6M4zd9r1wpXpSE1V5mjfNE68n94mN6Nrm67Hoabt4vBzfHmXy1N
jut80AgqovX0zDasx0jIrzHUuXQD6RDI7O+vrwEGk+UGDGy8Mu8usm0wrOqQ9fP4
QHQxYWZR+WAiGycXrf1pPNCVaw7bEuaCSyNf+rFnx1mMWzKkvFw1fM8VVO0oYsts
/CRxhS88tiE5edzajH+fJzmPDX+uLQTL/dgmxSD/BqwJ3f7WPi9pgmeCLeUN5R8v
RlJEl8rrWF+/RURZjdPqDpxdBrdEoNKwmEPkQHkPgJ2PHVzT5bo8AoYV3KUUl61r
EALQbr0mdDVXk16zswXiqZrkIi+5SMeQ4AfmuOkgg4bM+ZYIvqGic7JZVYwFQDwf
q/kP2bum7ASdumRUu/zg4qSPa5qwtvxbBpw27SDVz9t6n7g7ThyWcC8y6A9+UEVK
UP90a4iK4+GyomUw3Ou3dxDLbAnHbz9dfsPHGC16sv4TGyC4gKC1jf2s7Qx2sN8S
U2lzGWJhEJHylmXgHdliu1YQPRm4Wf6wvOY0Zg6FrAyUJZN+f0s+b4Ap/F9nz07C
zCTOyHnrXX8GpBfB23p6cEYFhHparqMXibSUDXpF3Zvnz3sxzou9iob8ZAOWyMiq
wkQuezORCR0uT9X45wmM7te4zhsGP606gP3uMTqZ/2MC7YlsC5LA9kg3tALevkzc
PSjpT28D4wdyj4v7+RaRd6fwpiFhju1ccrtspfcwXCkQyNcMr6zYv5cQh0C5aVbo
Dn1K43tOhisoPNKOWIfZ4KcM4vMNPUYzJgHh82cx1pHgCDXsal17FUJF47L7DCXc
w66srvL98K0MLcuM4F13RiMtv9o2dLwer2O1QHFs+Jwle9Kd+FsnRDVg/A9xHJnu
VCZdD/166gaJVpn/roQn6EIJJ2qFyCbI0kEUl33DvL5r1TQPPF1xTidPRukyBaxV
SGTssa6jpFkNV9j0n5HYhSL/an6SVhxb8UsvNkx642dKbRU14J00XqQE0c6bDrQV
tBJ84WSpdZ4UOhGe81qj49mpE0w4scRfeB/AVJwuW+OexZSMzLMTQKANS/RBQCNi
AFV8JV0wkcuiZGHZd9ZFhYvbW42x4G2d/R/W2crXhfmP1MR1ntuYxFxvsJr5Yy8g
rkz4e2fT8gfYmsJYbo9z1Pnf3O5Y/8lDyi7NCRzI4+EkbHQkht83mYeANp1wD8Ot
l8kRTpjgmaHuGDsML19RsucbRrggORbuJK4trgpzTU34NNG9uLEJ3g1d6UuW51A2
MP/HVy2vaHOUDnbe+LAIaMGXiixAT2bWof15eX2//Bdekb33LozPwr4OJ3s9EK4V
169uJ/t2aJ0UY8ZEWw2t7Lcr6Z1g38n8aWmFYIvEY/1yRsDAgNVAttj5GZBKb81i
YDGcqi+HBzSjmDYxH0RNCZkR+dlb/rKZPQR61/0w2+2otIgsIVNBL31tE6JJNFZS
YgdxGqXLzsxP1heJj+plOpYtwe3DvH4qecw3Ya6cckY2DPEjeFibMQfDABMKb4K5
M84DwI4CaOOIHI+91PH+FB2jUzPjN1i6+ukdHfrmtw4QkDYe8HfIyHJ4AzLAAoxe
FjU8v8eDBr0HVkZqNZZjKoRXpHVQZfiO8/0hTw4sJahq7NmymRC+iLo7WA57DAiS
/98mjTj4jSCbJLsqIKuG+RzQBB7sZHwqCXrWLTTE6QjZUh1LbSzy13sPrJmStiVp
gXgFFjPB7m9D5/hh8zyQD2gMLjHUyvQy4s6AhV8HdZC0XdcilWKr8UpG8U/tQxgM
8EDyi4l3jVfGPyppI13IAWZZTx3EYMMI7st5UXsoEsxcePvwSzZzNfKIfi3oYpO/
6bNsb1PcmGNZBSYuHHfd0K1sng4ssdJwnnFutOxCk1QX9f6Y7g9tnqzTymMVapPK
YduevukkExdnhhztlTDnm8990hX/vdZYCUtvP/8EixtNiOkzZpyHZjEewIx2hQkE
IUYRknx1E1xcqPgAe8hpSJt7/E6n0od5j+TuWoV0T9JP3V2OQ8IJnLR239x1TDG1
b89B5NzaxESYb3KdRubo6aTEwbSaA+w7dsk8N3F1l0mRuEDoAzgrq2x3UZMMweuk
HoXLakAKGoFF26WOyCx8ktgn+U06ZhCfDvGXj4kMeJ8tQCnORwDAzWTb2SOF5Eh+
zV/wBs+7zfX13KSr4hiNL2GgV96r2E7ZMZVgDFRClPqyrtJVrgfgNsgrbkxWSil3
Mv2t1q1sYi5eFdZnkFJdedmC6ikyD2jL7t0SAnPfACGxCHnjgF4wWY03sj1O7i+O
hDcjc1Q9/aGwdjhmL4ULTX4AvojtyFfasoDlbk93MHF3n7Rr84uCJzuw+aAHgJuE
szGzbNIG05DHFucxg0wBCPoCqrLvKYgVFeqJpvJ+5DxDoG3//2t/eVP0g3MxNxVq
aT1PdqWv9CWZfSwzPSF1zHIUtweT4hOW67FkGx6z46k1+jLVE6wSZh34Syc6s+jp
C5qnHNsBMqnUL4BP/tU6Z+5g/Of92p2ERIF3PcLWDAKi2Lko+HKqkSLMXPeQC6vf
7QCC3wcaEzHljtVCESyR+RBbSksxH6VUP5B5qlmzbi1l+e03CdBkNXtOD+wIjTxv
YxqwulkmRYMbCP9bmotbhFY+V/JhfkWKoplZglKvMpgY4UumYXEITR+onNnkrC2E
VsnKX9kJTlYqDoq9plhle/PulpCF2gKYVDkXwXRYNyIg77+g6YVFm5rDutfeJPz7
RdBhfv69p1J0mmiM20sl6qe4dgYuPk9dTZGoevFL0GEm2zBf7Jdxl/AENKcsyWYN
nPPRs0r6G/avxqbWjESFEUbfG84GT2tWqYYcEV0OBiVJaoCsL1+QsREKw1Ir4sf6
BYGoaTmbM3wC1rB8B22LBC7l6tiJTD3CA01u92RWBVbqalo8fQu5i5PkFqB4se/U
W0+xHXzrXU5spHeDeio/GW6Ntqj/fgzdYDDVz4dsjFHbuQVk29+KY+ZofLzm/gWq
GYxp6aVy15vOfKWNjLtxjCVBufVvxfN1QVmgmfhnj20k2yHD9GV3OWAvBdkEGkkg
f32gA5SBE/v2z7WeOl2zuQqDR03o8NT440R+VRCSMMAguz76d72FeEjnGbZvpqfz
fYNwsQjpghVywZ1j2yKKb4p9PQElrWhHjF/0j5n3OS42cX9FA2N+0l1H25DEqzRu
yRhjk9MCzAzI1CmKRyAWTwk07LF+BVnuoBdn1kMVhRkW5hIYydmdMxk2iTqlTufn
I3ladb7i0eaGC8TtbrVqT2pdRdwaSgPp1O1mci4u4T4QFJyuPeN3DnxvdJI00WlM
SE4J3SNj39/YEeRkvK4I+/EwFiPFXenPnEFuiYfXCVGw2CUxcMIFeRDzhCArLGs4
SYHlQVlH5EHp36oxo6t8z7oCrpMTttnIsIqxm+p6oSz/fbyAfjALvqHjlnLTrZXl
Ha1hMFMA0Zte7l+ZgOhd1EerJKNsPaWQPNgtw2iIm/Oa6cwsfPQM64muw4ZHxexv
v6b915PuQ9g7dkOowM/7qaSL9uGunxL0vFpjtEXkbNElvuxHD54XgkOEe69oHMV+
eKALRrp1OXUDIyU2GBlnqhBMTjA1QZMrjAKIzYbOOXK4CSL14Rwj7MnDO4oxP4FH
WCZD7GuPBj7SU9Nw7hd9n5/om4b4vTs4laRGZzjnkdEGcuFvmPL/YjwHl+3jhBOE
YOm481O4blpSrr0lh7OsIcVp9HG14D90FMQCeDK7DfNnF3WkaCLhNMWbLW6H5SfY
gPCBH/FIW8ks+B8Jxs5gDyOfzdGMrdsIKII/lJNCyyhnsT9rHYKzo8ugygZnqWVG
uEg6Xd9wWPPBi8b8KgpxmXLU+30DkiREFEvv0OJwzls3iZy7FDDm/qwFIQASYMTK
BvhymU7JqP815MejK5L9GU4SjwFXkqqR6iwjQTMRbyr5wsqND/J/yRRagTUvw5NH
THTO3prJkjopCMd/io2O1GR/VzZNr5Tsn01RwuABKmNt0KktWNia0nk0mjVf9fhE
SCkg0iZptZHvRqVsuu/tUDhnbpGwmlcJ3sgufwO8zHj44k2jDVLj4reE//LPAV8c
sSL4An9KeeaMQI9qVrkSLEj0S6uRRRLfGZmz6DiMMevxPBBgfGzCy266DHMraNr7
YAq5g5lxOnAG1iHi9bwzWuW6TuDiSw9meDE0P4hQ3QcGE3siAdqeYLUCCC0YBw3q
vUhzfoisgrCYwJpGElOgiBDU0cUX1OzzpuX9m03BLgj8BcmD35WKYBwbc9JGN/QH
zAYWV8VRDOb76/qVCrvKUKTB7dvRDtADlejPi9hoGlOiZBYSY/BzrZWZgjMFruyy
WLkFfBMs/KcEOu8stGp5cJZD8gAr6bqhHE/8E9C1WbAx/3NQCaSs+thrAg3Cn9uV
l868Y26L25i383MG+vRuBGs458EXfUYL/BiSTB9udyfsab31CdSRoT20xEx+yGXo
89c1l5WC/D0xackhy6rlLpmL/RqOD4UdV8IBJsn6QQWswuOYW55rSPKEew8YHFWy
ld5kZln3klRCUFm3Mojr8i8NpbLiAu5znCCAqbNQoGZHzeFEs6/hrPUUx95XfbEQ
62D3Vhvf/rsWwGuIlUjBoqIroi41YJt7btEkkX6r8+lcX8xK3HFAnz1s/pLsvrX8
Bs6NNXL388oRpaUR8CnJRldlUWGuqHowJBymv8Tp08y1qf3Keu2IirgplD+c00Do
+rfvsPCUwpM06wP6ctA5sgCtND2JkyNrNwmNRdn8SWu4hChIqs5XW8buTfocTmon
HfsUwWkDMrihnScFYPHeZUr5NdPIxrVAqtvDaeyD+YBLBxjoaAGOs0kgaUIewUZK
FVASYtBCpECLmti7+AtTzNOrB+oF+gqJLrdE7AVXnn68nu4OrgY5XscjMPJZNm01
uqIkhHAZeFaK6mBSbEClDqzvw7i7ST9aHoa7pJBkanV+Kg3hRSEDlswJVl9wWPVk
rbj8Un9B5bxRXcJt34N6Z081H/GTYye4c9ko0NI0IEF5P/x9mpk5RAxkHK8V86xz
ehXACAZx+nqZkb0Z53g6Yr3DB9TKwknTlhXkJuZnIHCnf9XxalWIyvGwdnmwKsu3
UOhnz/+N/uGSZQ4RFN0CVc+oPCiIpTmaBB+lBe9ra7ghjDcp1rA26L4mZ2iho0NR
soOgIpREN1TmXBvdcgz4B+NvCaMGIyLef8hZsJHN3HxNKrfJZKw7B5RLhSllYHKY
2djKpv7aeAUofPzZHnilT1e3dk2Xct0mFZQXfDB7syCUEf5rYdxDFPiMrDHEk8yC
6pZmchJ1JSf6yg5AVnIBlQNvB7+BeHrfesPgt6/a71x71QoPwipjAcPDNPi8LjhN
lG1OaybyLfID9mJ9gTOPKOO0gbnOdWM2AoayNpJR1DXDGZMBl1+8AwksS3fLD5dH
asmI5TpCJWsHElqh0SLgCRm0CFb5qFjXDcbPcG3l46Hgz95gmvHRYXVaIjmh3ziJ
FeFBb9usX7B+RenrcYbiIDj3berSdAoWPIccYRNRQ/DJJrmcW7dEWg3VUam23och
kiDeEqalJKPoi9a6nPdPR27XM7k3Aw/XnP+iNJ91VH7i5ae5f99c6oALHpbjj/EX
/P5qdcXsCngMXhVbqrUegRPeMwlxp0ClGsUo/uYjKhQHHn3uQ0AdPC2gF3D3hYcH
wuyovRXFA08MpOTJR0AUu6OkB/0vshY/r0y+fiIh6sxXzTjJ0cg+RsUfhN8nnEoA
boLmSZjVoF0ICtm31LDHiK4GNYWCHAFyplNs5SjXrvAVVaD0bcGk24G14Q4aRz6v
8m7CUJu2TqcWZbcLrRt6kxPbjXUTtMpTA0cYC6VPJ/Fe4btbXuQtGrT6MAIbS0HM
KgdJLW27cf6gEsMGoXOolFi9hX3JNXxEQbfoRHVGkhcaIsneq12Z77opKDAtGsKS
e1Hp2eP6oKvx9fOiD9WT5qGI9itaB7WZm7JeSwEyWpjKJYZpTErMjoBqrabrA62K
Wyr0ChCCkftLZqeReXP3rmDm2XLxexJH9gMRP8nFX+ua2Qz8mFDJWmVX/fjG7NBr
KL5UdYfgEQISdmG58zUAGNEu+I0xOXYcNKkhIQaZo0en26aFBj34qp93wNZcHHgI
TZyNrWzHhmSlOU7XxIXWxZgObxEdjYzet8DYohSYGhLNlGG9vS/8mxa1jiWyPVNY
gTcGxZpPkllUindy6ntqikv4G9vod/oGULEkqxMJBZUCiI850sPwsi/oEMgpqqG3
tzkB8EhPs+OdjgxJRLZGbVViIz6mOjcX2DStCtNxAYVujiVwLoAWEsYi3STCeupo
8xFLI/gZeWuFcHOqe9MopIXAxcCAEv04t4O1oke8lZSWnM7RWlmuQa15jt59/UI+
5fHJ2U85MJZUR4pmmSapUWFCljYlLGCyOF+iECjjeS31Rvgn+a57g+UUKJ4+SQvi
RBTK+qnKSn0NOJS/Gj5HfT3DL1+LBvZCLjCKp/fhiTSHQxWAaho3Fu8AHOKD3Iit
5lJQvhx6DgLMmF69B7K3GwjIjAgMi501dX8/ZXHbwGPgEPnDBAhLeTmYXGLHWzTt
tCUR7t2HaY6mf9w7TJCLFdXP3NR7GZ9TSXdz76FftCzF8ruRc94Ge1ckLm+2y6Ng
7EkSB6p4CDbHS34JAudA+LXJF9wP2xf4E/rLjB518RxVjB51mssdDR9t9bXXY7oG
6Wmsa+upvWJP91sIYbO8aA7BPFW/XZJ8Kq5GIM+5iogb9cAl+M1ZCzeWoXexgO+p
S9QsQzppM3v3oVfRQIXPgQhFH6/p1opon6XASHfDsLDHVlrhkhtfelUWNFsAdvgO
PpQy2bhvYUYnqq6+1yhqwa/nd4/Ys45IJZ5KLF9NyeWI/Vaj7NknUm/DQrsBk14U
0KKOD7rJ3sorxKaSw1uqLLRRF59PQ5sEZB75Bfxcq6Ai6kKQ9jiWWjnV0KbySn5f
vAGxVA6iiu1drdn7/XeahRUbQC1OnXDKtZSpgFj4DFkoEgfaefFCYVwBsJakYlhn
EZjwdUzJXL1ls9TFyTDU0oAb7DMOZDyI40zR9IWZfZA8VrUm6GCgnqno6S24+Q0Q
4/FfyG+Y79bA4ibO5wk/uo29o69PBBbcJBb5Ci53CoFJImbRCysnDBSK+BogJwNs
gTMUfgRR/esuN2kdLOnJECS/I9Bsy4XkXORCoWExvzRCj66qKfQ3HYVZWdqEZa5U
p/Btl0lQt9yxGB56ESawlZ8MNEXKwG/2rq6sV6nQUUp1uO4EJA6voLwcxkNtYFH6
2dkfRe3R0ngKQT+wzQN3MRYhFAaCO8DOAwO5rhxhivEqSuQBJt6Al08oDYc3OBjr
Pt+9pmE7b+lCb50Nx17D6whc3qwoFEqcVea5OCdzGmmZm3YVFnA8QmQmTO3mmVdM
yDNj2IwoopAbAs91iKKtIobSw2cipZBPEA07A6QD9rbtcvzxFnm6GllZpctdM2Cr
SLTnKOF5K0uHwvPb6nk4TSXnjw+hrL9Fw6eDt7DWSJmsiH4dZYcHYOhGQEoSSFGi
o124leejYn+MVGYpV9fHXYK5XOHxBDT+uv1ixgC6FTvvmP2IHYtadYyApzgUa9VH
eWdzMHh2hz1dHUuQ2Wym7iutEnC8Yh5Eio1jI5EG6K0II/pgHrLTGN6LTq60QQ2P
6P/CIeugP+V/pfeXwHlys07FDdDQitI0VrfoQBmRqpVnfyBFqK1+/gwox5n6WL/c
HOtBj1IM1sakGakQydzWOEMkutUV0qZjAAacULuvw+BJFkc6my/50GXLYZLw+4Hw
yQOM0ofCNYX+MWcM9ysgODDg+omeefAe74dyacSpURtUjF3zi87GYh9yNcn+WLlB
prGZk8Glp/4P3OMpUAdtOrVuplP4xPsJ45mnL6WARf8jdx7bDYuUdOVGWV6tq93z
wcqQkZvEhPcskqgZO8OMCoDtRfKdbUEPd5fkTlO2quLBPV3WYNDvl7Mwj1Q988Wt
6ge/rV+YAZ2+orekXlb6EBDmynCSXcKD+WYLd73DJj6inOLvNl5FE+5SL0ZbU3Mr
5u4sX0R1tTPJn8yIGL2PLIOUBuq5AAlYLUCnibLlg30pCVMf68cUDDdyP1zWjZoX
AUpDBKWC+5T3CBF2eyXKKWQ8BFFJMaIZE8DLPprgVhuDqkeRJJMNRaSTQj1jc3KC
TuKVAXvFR70DNsGGA3+aqa/U4OXJJh1sxCeaoj0risKPmL/jOLPGnZ+XSFwv6Ren
XT/Pb5nI+JiHIzB+PN1DbFvitbRQY7PEKmfOaRv/uYr5RMR0rnCQLrbBDy/exVLR
4K2lEX6H56TlfmgbbsRZwB7/mpJXHnctMkzJs8PG4VmiNeGIoNTGWDhYhqqKpmCR
KNn0jjuWny9UkuuFcS9iDk/RUk69Kyr3S+RZPKzJU20W+DVNKMLiUktecR2+FMlN
5N8nXjHoiW6FALhBF9JK0Z9RWSiVdM80ia1CeS8lx/0FJ0iUhNzb33VNDhf20pXW
oQHXzWs5bcbBzVu+HePeiCieHVFCE5Vs0mr6uFSVizbEIAR/OQ4rWArqpkunkAJF
5Rn6vgZXU4MZBra8TXU5Ndol2S7qB30Ac20PpKYt9iMFhNYlncS/SBcVlBqIqeO0
0jLZQ780AtOSelzYwZzQkH5r16VZobeIrF8N70NXFnRjBP5eWhk44L7uyLX0QpzO
aGcixBr+11f5/wwEJOb64RZx1nTlat3B073i04txq1AbaltQkvnLHEMGdId2/svY
ZZlG2UILUtouMPlU+mOwPwAQrXKOeLvf5COGhJnt5KSgX3C3v7S8DaIGbr3OTU/5
pRnsCrjet4yGJx9K7mNgKofqJGqLSMwY0u8WeJJt4k6uCE9R2H7BdfFVU0p0Xdd6
pECtjmfKrpgNgGmA8D32KUswK1NMeUBW+v8F5UlX9G+v8NaPqCEpzmMFnetrO9H7
y5z/V8F1xnlrAgbl9Z3rW2WOUS8uX1UxN4gXCs2E/Z+zNkGUDWc0zpQP+6qz1Q0t
z+VZajckEyq55svDtYVYbFdomyTN4erXAsfA1VOZHAKXyLrCEMJsoylg2jKIkOlB
bhu/XlbxOAwlEU7m+v6H5/jR3A8QQi9/8MSb+KPLv7O4RRmYwcaEz7fK/iJK9NQB
msrUXktGNvKH/CO8EjLIsFUe9yBVKYOEimkjWMjTyD2fzoLUcbBxCV+0OSlh4aSK
53GbvPfRAVGJDGFPvMA25tMU6kpaAk4cK2MUjpzNaBnEsjE4Fk6JyJDVOiPN43+g
gX2B0qCulBHNwcOcWJ8mBqU5YwhVHDSGICNGPgQ/XFK+mf/eMV5TqEdhmMx7KvVl
bSDaKNL2NSInF9ZA9yqckoeCyrBwt+5+Xzoe/3w2Sdi82rzKDAwYlGewIeuPhjYq
5bZyv/A/gi9sdim19FuSljpGAsmNp1ZE4t5ssxQhr+ubaYZfKNBhOvs0RaQAKILZ
08vDW9vVtoMw0L+kQWtr74SXpG0nRhAPcWV8bOWIXeFlpHl6mPfIWCc3HtI7kKil
3/q+hpia6MKbuZdas4dV5gu0nQ1Y9Ta0musmD1vZsF6AZen8E77HoVj4NAWvWC6i
j8/c7i2niIw+rHk3osTxmhjRz6pUZ42kO6YNg/P66I77JG2KmL75vRlVvvTjZ3VF
aEYjm7eip7l0ut3U4tdflnkudEvM7rh6gg6EOHVh1x/0YiloWgfrr8Qat9v5x2Vz
eibxoB8rzkP2jTN0a7QSX+CxnB2389sJ/LTtglWDsJwmcXv5t+/xXUChZoky7xre
gVWyQJ2dkXy3KDe9MITKwO9LBZsDUk/leF1/hcrRUk37LGx0R+P/QIaAQTTggx7z
89yIt0H+11vYnPE591dI5AWKYAF0PXtbwCJcLNGY7T/CL8bDgFrqDz84zDVVXzus
IiRFLs1mvLg9SDe/Ml73mg4zlDaMeMXnN+2cPs5tRqSQ9g9KP/jsTDpd9Tx2qmP0
uo5gdPQcXX5al6nRjD++h+Ri9dfqZ9EWx+q1ExXw0GNgordNzDd+YP4kdCVmdJIt
W2W3aQh3EQ5eUYU84piboNbXedxRHrTC2EhYATSETw9XGt9fb2WB8/26TsN/UM+G
KvQNO1ULu4sQ/NOlvA+pBUoEZiRfSIKGAPd4w6ZuFiY8wL28gQRID2DhKyUkvoO5
Ivg70WsB5bOeoDQMysy7CjOZBXF7rjZI8fKqRP7Vw3omJlzX4E2iqHVekRTHtZC0
8nMkygCo5ecg5PRaVPp/4ZCboybv/LDkdp3acixng4t/TG3Ohk4tdg+2y6gDFhvJ
nETB9Jie4N/NsBmPgXl0hq9omwcnVEh6ifTG0Atb4id2kCvfKq033NHLvdjF6oYb
QCbm1gWMQm+9JomursNMRrvEnTrA8EqtmqKk8vcf0jjh5ODZK2AoDL02WQlKtvKh
KZoiAxGR0oUfp5aFNl3+vQ/0mERokV4RS9jSeukDUQvxsoU1cYea3b1XMnWxFRrw
3JBDCXDq6mkP4FKbBQduzItWmxW3R8LweEjmRhbCWptgUSWb614cXT8QGAs2gEJ7
EObwc/jRBm7wbVUU+ywf5/fVpHvVCGLYtslBc2q0NYVjTjYdckJJi0DG1AVbzqJw
o8MDKKxL8aQa0f6mHZdB5dtbA+3x2YumNYt+Vdrkn0/p8jhEE1GIja3uK7+CAybN
658IKKJ5GVVN3S62qYVru0rkWAJ2HN6nxgu7oA7XbIvGzstHHlS1kvtLUYVW9G2H
GxXIi5ukwZkblSDLNrelenWeoFIVG/ahl8ackodhfZF2rjJoX9OQMllh/TBq8jOF
DBL6OajjNS5c5ViIJlbTxjMWsTCmcsUyfh+ko5NvA3uqHs4NAqQybbSVS0V8Tf5Y
Q5ZxQhruZMGxkRX+Y8rzMt98NLOtIrTdDm9BgPQ12z9PJ8wU1s7GJjETs0SG6xDs
hrz5ZE0KPufM7DP5eGpKlwuthxbrnv5VpQ6QlnCZ3IKUQzshCsx8gBz259VYWrGW
C+uYV4yRvrYxukJRyOaSY02cp3KwptDEmTn/won9P4syGrct4JKN5YgvWxP32Pqh
e68Px1vjNkbcfEtfCI9Za4Fu7WLqEOVR5RuDUiP9DL3Tac+OM8GV157e/JLAiFhQ
OK6GNwXE9GSQYfaCMitutG4vcOZwbF8iqpW2UKk4JZskq/u8ID14v65z33ZvBk5v
xeEoHjW/r0uUp29iPpvKnO94eeFWYBf6hJRsewbOXDCcOxwbIvWdqmq05AM4e58A
POiQ54UOJDkpyMQyqSKvM4Og1AHShCvtjJR0+r15EAgDg1uZ6TVTP5+FA3AjfDjR
QSn242Xf1X5sGe92mIK/TmPUj+GmMpY61kFAgkyPe4m6zjx6B/Caop4q4GbPK497
nbiHfdvb3RbU8YgiXBcB2KTeTum4Tl2FgeVVj/jQPZm+Ul4YMhzaIt0H4TpQeDe1
E6wnj4+M9wzbXzGYU+3/2XbjKuOQaRA5mVkjml2rUgQGbhpf2DsesNojes5hTeKk
F9qdq81cIBtuX4xJlEJabl2H4eAliNB6q5D6VAo6Sh1d0ZwHOA1PKsBEsbJqfDb3
G4k/XsUTsyU3vMeuNwyRToEs74XjadU+fijak001donE/YSs1pUE+Pl5vnkHA/U9
NMI4pjXDKI380V5xE2ZV8w/MPZ1tl4ejlUV0Kz/WSkYsFEHoj/dEOJUb6v2iqKM+
z2etEps2EI2eiWVPQG7n9loZDbrhFah2kti+10jK0AfU9n15s6d1BCt9HRSL4TXy
av3EEqIeqgRghLIU89J2sap6T3w/1XzgWRbskzXvtp/VW4Lj/XtsnzBI0cLRx33w
J7yQO7LOKAPSVGuf9yhX7ay1SZBw6z1HsjqD2XBmDy1kIJ6A9IAKpQfUOUPPSTRk
hP7wKUVoQmg+1Jnjl7F+fUV/fRRNhGT8ZBwUpvm1RrynbwgVepz7Hh786zAsEv16
93kWCcuoolRR5/bShI79zXQ1uupFuX1pokFxjapL+xk3JgOxGWN/KqMP/THtx6mx
yrryzreGz0JictqF8ZxanYf4MhKUubWMvxLe7GanE7RzdPuXBUTW5JFQEM3JZaUM
ETPoBD83J9meilXh09zOAXLm0CQUu4eH2AdZ3MlX8YJApy8ydl8sUjI0785OyhcW
+EBDHgyIbkZ8rJILzlns7I2Lq61B0QoHzjB99xwqydRqAAFcY5u+/lNw/R1tAfMA
33ecfwgzgOLb9v+2JOizsj3LbwBM1B/JZG0ryYPdIkv4ztZKKWtXSFiEs74mxEd0
cLZuLOUQdJS9rKXlMhQ1iRHLqmpMOCT9OM6EtYwL7nzsK78mb+H2wP5EzlKbygJm
XBW020L4yxTAjR5zmb64zQLkcz0GRhBkPm64UfjYiB2ipkDVyQRpgsi8VeDyx4ta
fN+VbxRDlqDh41JyjiTbFk9ybYRqy9y1uKXRIXilvqlf9HvzHcG1/bsASyyBHH/7
Q5w6oJukuU+6a2LrO74UFHxMlaUo9By8dGFdp7LmDBs3kxGPdgPh4t8AQ23jm256
NU90inGinYRkk6958I7lkL3sb0MPDujj4dkWFs8hIIFuvPngcHmwAgFEVG/PdWRx
oEL4XzHiARwzJOTyVo3n+P5KLzucbkvGNj+XM8zEMbCW2taiIIH8tUg1u1UgxBHV
ir/AU4LqMcfIVTzHHB/POs3DUqN8pSyVL9mtHggf9tUNa4EyYfIrvrOeNIsw83CE
nQfSjuCnfaCYHUBuDe9prucvVD+PM/vg87j3QQLYOX8K0AqZVbVyYfp6o22RxZk5
tRRuP9P29/7xiH/+/wfpdQQC74xOddAPMjkceT7fxlWWjyFdzshPtekzg93+Jy/o
LJ25i7xeqrbpst6D7BZ1vVN0sM740oFyLxpPUhjSj3TaCqIQIUMOr4ycM4J6IbNl
a0qImxT/cwxB/xkEU451MpNvRezKlxMDAt20KvrCvxsmfEqgdBWKYvU6Z6x83dxn
WORnEaPzjaR2v202nf9P/Mm+X75B0pppuPa79r3ZDED2VhUEWemM4+5CUuHzIcbR
takDd1fep+0jFRLEJXmwa5Qcl3F4wld1DQ4po1Zzl94PPZi8ieZrLdS36OM4H8VI
M2nPzcZVIiM+HkUjWmix8T1MIf7TqYn2fDp1baoh1dMN8rw9P3xaX+1ZLP2y3DAl
mProWS93F4pk59xt65BGXdM8rcu73qRNAjf0Eot8ZnM566CcijanND8e2ADW9fK4
DGugqmRaq34KQLjL5FWIp2JD8Ef1DuacCuOBi3shTERF8trjgUoAJdHgyh7qRf7M
Hn7R5if+E4hOXhNa02wxQTfDerltJ0Qyf/pqIDjFzhzy1nbtKPPcHB+Fbrd1m2Hv
XEhyqU7zqEXTw+g+dmkSBrIj4FUsi0oUqi61dsT1zmo8Ad/lh2+LNCSAbXyfH5+3
Ipq9FkQdmlmRPcqwlJ3YrlAjhDtVpmYwnvh5Hzf7yaO+BgBR1NXLVUOxPLVuI8yj
AknegN+yT4WS0s7DE32tBM/cwsAyqTsGInVM3MDnEFD8k/0QUd24dwSL8XQHRFaa
O1wo7qL6pD2/HBqGUmfnBR1zT/9FFR0r+bEo13EFE+PejxyY2KJ9GQayB/9O8reI
RYqmJ+iSmYitEe4O/ZxRev2J81onwDd03T9/QU7TH1VyCoJVfGCxXZO0wUzZOnly
Q87Ud1FR5UE04oDIDg8In9Jp3C3OUK5uMIkxuhirD4Xgi5weqlTGwWVz5e6VSkA0
+mhA8pKmrf+CE/YROEEvS/xXfk2VQ1Jvun9gPSQre/+Bi8P/r4BQ5MLjY0LRGFH7
6JYdr/O8JKKqvQkSHaJlmPcbTQUmFgyNEzNx9y3rjUrZmoBNPLyGf1xmsRs1JYsq
vDeAOTARYzKl5vdXscnTlIV3rqOM566znlvqcNh0h+St2gW2Np/Grdan1/akLu3Z
jEm3rx4f9EWLqOCW9Pqvw/+0DPky55yq/FypEgULtEk9zWbCYRvh6MqHdm4b2oe0
rlxKUPHtQjwilhgmcGGavE0lJxqTRq3yQhmKt5La1bZyjNU5rK7xQqNA9JgD3D1p
qpg1o1751uridNF+PTqPYFsnMpXh4jVrwQjDIUZHrBeUKen/N2ahQx4qp7ZKwNrU
OCC1rLMCFHW6HfA3lk9ZFDByps3Kw2zyuJBPdNFxYAD0hC+JSPPjZ9i5CgQEQDBh
OL+Uniby5ROgvwpbbv0xzrIIJpwr8qu0XsIETWFfonIAELF3KUgoZcpE3y8Q0e4T
LxrcN+85uidY8baRaU0+szWee+uW90sLvT/CQpK8b47qqzDyvgTi0p/5WxjKeUJx
nOtF311yrWjP904JCfrA+k5hjV/VqJT8REy1uNXTTWNxNJddlvePxnNAwHLAcOn3
2Lk/PCQp8GcSDmp0NGUu89Yx0JwoaBRiIQANalkCfWyEbsfSDXTTFOdYW08NEui2
TaGFwPUIUYXtbxwsI6SZb1YoIgEUFARqzliQzk1NaAkHLVxKwSpmsvVKfzz/8uK2
odj9xVMSvYLUCgMdREk8W4v0SwYIOMmFy7TriQ4hCHPTDfs1J1SUjBJnzTsjzwrp
B97Eg0phTRyJvOptHPjF7lGy2bgI/ezNh7rGPdxfSrTwZpN4jG2uHXpHot7id1P6
BAmQv7YmUfqWOB7KAUm3etSejwh/JsYAeNO2oLyA8VLhJQMNhCyyRzSrQ3tYlc2c
8UXqtorFH/ToJiUchcPfo5oCPM15JgEqLVk7mKwVlMnIdqcPRBhd9dFKHW5Eyi8Z
FHM+LHPe310kLjOda0EMgu63I/Jtt896EyVwMESuzA0hgwGcV47CVa8n5Zg7CuIE
wkiV2YsMVGM/e2AJNyQU6bXGBhkXUVsjU7qYS0AXcUJOOHCq2EYiqmPXqI35ZoNf
I8E3CxV1XipEvCHZ6gujOK1PiUruVXuw08uPxRnq7aetxDSbGN5lER4eKa/rLFhl
vZzV3bebap/7MdDOAGqQ9PGUAELjzlfp0sjKPFEvCKQUNdsTRFyeKqGNu6lnmbvk
sB2Ogu20fUDoeLCKQMrkyh0RkAB/NER6UsfVRNJdW1qp1VRuIRSw60yZVNbfu+yK
0HujD0NQJasJedGL3/JLF2QrxpHDuGso8rOX7bf06EBUXFNcJqIoFT44AvH0wesK
M/8lK8cPh/m654JmH4RH/bI71chYbp3UsIqieBU86dRJr9tIe34vGOw4vZQCDENv
Gwj1cK/3Ueu6GOi/2Y3dtGA9nOb2Di69aIMVJqXTwSkvUuTUJ49fM9zb4Y4YW5yL
LftFZObSQWa3eUpzouhvY3QssRNDmYXA3LoMcHioC8R1AkveUNWg5kSHWHWLOGoL
9oop/9Qww58EP0UHLGehs61ObjcVnjmAEaEZj0zq6rS2WaIeqkvJf/YxbWbpnhWr
j8XdK0YBuJ0WFJC6Nb7Ls5yRTry+BrDHgoW0DASW2MzijyUbc6MleMYllzPf1Wnt
xB16aCA9OyQQm3JDbq/x5ALjgiosT4An64fgA3MVbjbc9cI6yE4ndzYjEmTK+A/K
NS9ZSosfIXXy4ncAN8Gyj4bZsc9LMzYlw1ueODzI/PobL+dHMi9FK8cWFufo+tXC
VJZXsFRGgjh/wLt2yDHE3E4EpwTv1fJzY1XVVq/Uzj6ddlsMaJfHKf4Wq5w2m/cO
2pZ0Umurn7bCn5r3WijXOGQWI0WyB1PY9Rbpe0eVdtYnc9gX5AkiaGVe0xRUYpY9
DdWSsRjAedAGOvBu3HXxOC9HivkH5VIcqc/jZSNaqQa0xr45Y/95ughwe1TC0nk7
rubbL7ha6BUNCoT84g8Y1HlM+IdjAfCX1ZX7y46h9orFs9+ntsuDc+7vSGJf1/PM
BMgbNhJHUnlrjyi6FqWcAFi2GKqW2ltp6PMy9WWHDX9WFa765dgpbsD+jnC6q9fl
+QsVKXXVVoHUvzCK0u8hZYTDFVlhAm3VShwNOHk4SKvEimU2cSHeoWU9SImsHgBR
jEL1OUcwVTIEg9O1aqzmgHPIOUdsXQuKd9cIdgL7F+47lIuZMVx9S00S7pcAQ7fM
SZibQ1rrNrlw0W/LasAOVBOPHf0rxff6MuM06uydo3q3q9eIIEdZ2mznfB/Ghr32
UYBs0TMl0B4ncod2Iaa0Z+scoGZT6+DpK/8lmY+8Cc7jbdR+goTgILm/a4363rRF
/4AE/Xn0p9/wPc9spa14axFyr5TZIry3oRqnNlkuH7vIJo25cagL4doqyzbC2Tml
SWkcPky1GUUfiJ6Lpw7keIRp4pf4i218hc9bAKknHaQfiE4CRYIg1cAx9EFa0Vvl
DDbYwJEmcZE7SeYyAowdkTmBb49pI4K2ERtUFN7Xf4Ic6vXXhL4HscQyjeEGe9xX
amluAFuEhhXUm9btLeGpFyK3Bbn1XLkhc90+UUcU2joDdQkgGMFO9V+O21BmeX2s
v8+BfTBDpUzpUAJVtgiI5ASftwRHQlPEYIfxYTh2BBQ1QDj9QWJM//vitduwv56D
GAXz8Ru3OPj51VaYeqWEhIY7c/trrg7lgo/Cti9RMmBndYs173aYkJ/hAUx+jmhF
JM+7/XE5VPzXJwgPlvSrUeLJPGafrSOrZWri2/meafH698w2mJkjz2P4viINxhw4
Aao08HAuHdUtXs6rSIJDXEoPm9RCvSY3Yvk436My0lUb06jRe9o+xusNcX1imDwD
osKOhpwPnu/p3bL5QZvUn9iuO41JQaEBpVH5BOAY0NGblbRlLgcbyXE01Jl/9ngU
i8Oj05ZFYpp1UA7TdXaoK9QclW574wg3KMrkhiSv89fkplwYPguYLIccSFj+Vqnn
kSHmfcgvRMd4mGWe3JEoUyp4TJBC1Fz4ZRB5MALIqwx2JRYYZxQvE2dEZxO+0CyP
IRNkXGhATzn9XhVUNb5B25HKVFGbIgXvZkQRDk5ISU+S5MSMp2E1qDGOmmZyxfnv
Bgqt0Nj4Pm08NGBdLd6ZNuRVdi5piStBUfdof3ypStj2XKo1QapsYTkGBawyejEs
pAsF09ymaXoEiIjrHKFoYpePeDwJlD6HDlrBAabewjGSD0cWBsO/iQelDazWduuL
o117gCg9bJgFFonE+/8BRX+w3i5zsTUPn1Cuaup2VrPSv64T12tByK4EeafSK3r3
jVOawvz5PF3NfooCe8i1sW9KlXAbYJVz5ntXomjPNoruB91Wuq7yKswXl6e+vq6V
kQm9QlAqrTDVieyHH4QLa8h+HIVxGfa6IMuLSm8Kl+LqseqIEcfntNXiL7jjqdQQ
rjSJxSZOfHRE58YOkiE04p6+grR9U30lSJjZxXy3D7o+B2Rzzz6MAC5rHC0yqEYh
nYruOB7YzDRTs7AfXu0P5dbItmqaiEGnHtTFC/ljZkDnM+o9sDYwYcyUExBCK/Nx
kdFX8lYJHq0Zt+KlC/WQV9gkpaY/l2M8vfU9XtoRT8B0KKd5HmXWJ1f7iz2mG7Q/
j0L0NT3bpxUno3M4MyG330bBDHFQAB7kDA0xMN42HbiWV8j941gXE4hxoplxNm44
payfu6GWPB5whdZVkvc9dGzmN5NnrOSweKKje7A27VFc0fuMnRTwKjDvTqf8YliR
JJB1eaoHAFLCYB/RuvdaVWG5DYuHXTC3rX/UMdCDjiWysg1uK4B75UxwD2QjZYog
Wc5LGP1N+Ch5XEkadHgDyTukKxRVEJBJzg3tNmGvsCPIGjQEoP7MaNvsKn3BgYFp
Dow1QWC+r8ci4zk2z0HeE+eKEKMEGJQ30QzZKKLZKeSDgXxcFY/+T6travvKwmih
NErizTEl7bfpMcVLuQj26+q4rGwxI+9xlN+yWo7yRnb2tQ/psfYegGNsD7BS44IQ
VQ9/mz4aVEs7wi+OhDEd8w9CLg9+NwV+3LpokUyFNwsAy+5s8vG0jH7tIivVvLuX
heXk4HCqvQapgAOz3BrRhltL3UDInEu9Fg1eVO6uLqHgVkC4eWFdDwF571Y9qYUY
f/961k/1HrU2EcoplfIhnK4aN19qbthhEUJXPh341xHlIwuWP+/E0FiOTFN03bTf
pcpGXHst5dfzUasQbuTZbvv/qGRLKrRBZkfyRbnx+0w6ZkLVwqdwz8P9uuN99LGR
uJzBmwB50F2ynYeyQqnH2Z+7kMXQd7Xz9uX9y0LWNtpHhvOSYhSUUMNpUuFYjpjx
XWqY/4mhSbgexwSC8ProsQ0+9QfXDdNbUdUSFS92pKaVHHwDJkRjubWM0EbHj5UJ
PJ+MYlz19hO+jIvRban+6Z3p8H1mxAXrKi4zf9uvEt7DLEtDqB2mcCjjUnp2FGFy
seOdMVYa6rzyOLEJzcR1lMh6NgjmAuFSlG8npBKovFPr5R/NxFIR3Ves3Sbmz0a6
TZLHv1gjE8rlqKV6mkQPquxsZHA1ges7c0PKo+k7P3CtgAnZxbQ41Njk/jtZYo/5
lJBng3AwuNfe8BLRuVRwQPwmueGN2alX8w09rHPZwKelcwTU5Ja/y3+/6h4sfzxO
xL51RXG+BSGJX6PZj3xL+XG+idsiVI9HNaBHNM8mtQKOzzfKXTAngHhOhZq7bryT
ydxKhAgaA0qDJzAJnHpgFyacLJrjuatTzqcuawN5Fz38UpSh832wYy0nYuBfeBB6
SE0luM8gEgJQZNGwGrFXyzZEg3JOPYOWjbcmUGVCjSP2jvnSTAF+g9gAkxjZ3E6w
YJ3k68tMv8prPDMfJnfW/adHehTZfEi8NbVi6M0yM7/YJszteHBCiJV9wLI8LHbF
ui0TJ5lUgeyyyJX9pVhIjY2oLqcR9GZ/SEoIGXl444UlsQa73eA52R5dEJ5BD92q
2gCnFIv+TDzY6CfDC5rig6BWrvJdQlxUT25H4KyDcVdhGPlVIAN1PgcXwdE0lAe8
jUuOWw5TNyAF2gx01+Ciy3c/cMFmb3KhncS/dmHId3pb3Zynytwz41g/BIbNNsHF
5uzcUnC70UJ1/XPItokpvXjKBcMtP/ZQkbFIx0KQ1scu63XxJa4XWqUZV1U0NFnl
jlYj+mEMAVxaEt1nqcNghFh1KOqHnOPgFyFIEB/uWI35HVWacOUmL36Snin9HNu0
anTf8iLedvhYN7ShcTSMS3MGMWthfbKwvYdkwaGY5FIHFxYgaKylxJG1Ku5rQ8v9
JQQ5l/GQdDyI1LoeK4pPbbA0NBBcHegwvm3eMslRj1B9yclKNCHtLF65uJL0Qwtp
oChLKIJKG6RGcWJ+EP+E01EHo4i+MAbn4k19Y5d6rcsbWM2V6DP/eV9x541kC7yx
ZuK+xKCvhvG5HiFtBDvDbwosPe3SERaWLSQxt7F60wOjrjPZMzvc9x14IcgCpqN/
6imXdAd0D5zdY+B42vw6FofK9EAbQ5SYhxqv8BuHlPtDKaXapw3BhCNH3Y6lGbhV
bqHrqktBShKOPAQ77rx77UcvUKd/Dqy9khfWwRbKSU33L7bWxVMdXs5DfsxZ5yRq
by8yuB/uHPJEVnbSn6PK1rgMqIQuT2eK2imxagYTU1VVwJRM/54XaMpQJFnnvqCU
rDxfFJbvFJtPd5tcPmZMi/PNuZPHNLo4hYVpwfftcSVxGBeNIE6No3ncOaMWndKR
V3mLFAF15YhwIcwmV315ANTw1Yc0mXkBEHdUkuN5HYbAVbP5vuakwj9r/sZF7igz
a1wafxm56GPQyjiJU/5htT57KPdbH7Qh5o2g7VHE3OqtiVOM1j/lqYF13BvWStl0
OqtqYTN9b8etz7Yj1czErkFUTd2omWKSePsBcfQTM0AasMMeLbvMmpDl8UNrHp21
x2n4JoG4HvH3zjn5IZRpZsiOprbvvwb8yaIAX1xIYe42WyTT0KSRJ+JYjWWr27wG
KKjwL3oQ5+rWd3TaBxCLSvbcF37gGUsU9aD+gCTT46VZqJjM6VWzkbDHcRAmfu3h
DJCGFzCtHq7kYoye3TWKWBUBFUoPO1dV6yGCKLoD7QWET3LF9oPRuYLQ15u1vFgL
wW6RcjPfrohktkCx1chdN+CPDIr2t5truF3fcNR507la+IXYV4WgzBV2tvxOHBtn
/19OeNM+UvuZZTKIG+trn+Sdbd7TEFGmaxhfySeB3fDmNiw8My64YMftso2ONrkL
d+a6IMseOxoYKS9YKof8bJsE6J6AEaBou4zmP6LOtr1TNOk/yitcRkwIuPV0HuUW
oKsY04VyipJg3uRhnm33vbtR/4mPFUVMOrk7iHkdix/FxvgH/iOSNdc3tjIUaMPN
5HY0HX9tZ4/gHNH3d0OZEH+Si+19oQbu+CNYo8c1e4o/YhKAKwTLjktWEe79dx6T
+plWEWI8+k2bpmWmymdzCiIH/15lOW7+hHmMPY/LXYTAyOkcrV3R1PaDGemztT6H
dmyLLQBakqzVbyvOHGiCIY0zRIAWGiKiPo4P6j5AHUXA+/8Z6ROucPTAt0oLnpkg
e2FJi39NwpbaI2i8YcP1pwT1vb09pPQGriyI8DsTgcwWZ4wtGiKrdzv8HRGoyEO3
Rb89o0fX0mU0mM4DvWeAJfMOZ4iiyKYvsjN8SyPxI3LPz+k+bTu8DbHyX2qNz8Rp
J7Yhydp62URsWguf6Bwwec9TqNrsJuhXy5InJCzNd5ATORxgEK/Zv9vLypsGdPrF
sSbBk8VraMLRAMU6Ud8M7r4XOIGAb5mq1K4HHID4LSVVTu83sWSJXboFHEV7RJBI
d+tM4HFW8sC9PPFwVWYHdXOqGKSBBBIeMT8qs4fftaOgKOzt15vCypR+SIsmGIJp
Ecc7ymDyHpPP1WVbaAM52c/SeFZv/F4lTuC7mqo/F51znSj4Lb3s9QKHLCibJvTT
J0gOvjArFDPl8AI+qkS6WVa2oXOpw7WZTW3U8SrYmD11EOxSsTYs6gA54n6fBRPJ
jYu2A/bqqI0GIUueRuwJ7TbKhCc4NUjGTVQtZVhZFvA7FJ0AY3gZ+8d0p5SSOFXl
8J4CK2n6hNMWzFHfuzq+2zdjMH1ZrtpW8Nw+Y6radmxpC1ttWshkKker2ayxXlL+
CpeKOAkSsXmZXPPsCtW9QELjUhpRRn6OnUxxQz6saQqKkcCVdmtmUbUs7rpCfuGm
B8Cg0T28J62T4wna0B8TJgPrT5I5ruoHoPnLmZLyo1JRDF0p3LuVELtO2hu2E8aQ
xf3OARA+knXDOK4YgOKxhaOBnvzjTLdzGsIC6ZMDYcETUYCevmcUYPBY8Rg7814E
k8nt1Mlt/7XemsU9yx/xX4nMrJ/1a6FqQZcl/8tOp0M09axB9FlmkNfmYoOqIdTD
2V1dcakiGfY3HdlygUWq4gx8eIMO/aS2FiE3OPnK/p1WcthD9V4frTN3BNe+N7Ne
31pzmfbo7zEGT45RJhAF22XPipP1LLzCArH2f59eu8K5EVsMgL8B2Z9fyK874d1N
DHuXXJ+M9t2sK6i+PcJXsM6PtYpkijwuWDKtzBxexRWALamFwDQpxZqDPIB8Y5cj
udMZMRHP2Ln007IR8zC/KrRYJBu6K/WXkchNb00NOsJNSZmbJ5WITmiMP1AFQQCJ
tae0oDqWhZJV/bODSVb7M+M/0Z3FdYvGlrwsNwm13qQtb8VsEFkUu8XKGOHQANQa
3V2kUFJPB2Nust8LCyZxa+FU14Fymqk4At2srv/f3pqCSZANY6lXvgSc8HnQXoqG
mL6plpjBMQGWZWCTUuo8UA3yMr0nx+XuEfm4Enwly9nA5L2EJElpJptMdZg6q9U/
VS04BqgEFyQ/XEaEWnQbhs7IS3DZoeaPHT4HD+RlHYj7KziAvXx4QC7clsyTy37u
D+bWEIqFcP0tzKkn6kMiOdiqpRnQR0hpKD4eiPxKGYyIfPgrJKuvClEFyNByIJmS
lOMSTLzfsLiSVxGYXurGAj1epd5Etm+k3kj9ctd3OsXMrMPb0bL5udMBA0iTs/Ml
EXrnvPAnUSumWPEcVqW9gEE3SKKf3dgRGkqh2dGxF4j0sBGNPL3US2wCu3NYAPvJ
34By+q4ihd/+6dJYamTLWjQ8fxHTKn6+rdmFg/mGGH3Vv0j+f95iDvRJ54rcwQg5
01nKskArHwndAM8nhmpfcbfqRjAYQ3Tpud+Xk8BwbCd2IrwTvHBRdPhTadoMywfu
6Ycm8v9rioaGmCmq7rc5j2Wj50c13MCzG1rw1lyg9apWDlMCKfIiukL3h/Fh+QyM
w4mfERXLpO/3+0D0LkO6FuscBsuBITiky5yEtk0joVL7y7H8VlRdN/+/MSnJKLQI
gz48Tc9tOsi7SCeNq8LU5Ui4a1QjgBGSDVWLo3aGn5vm5TRpG8X0r5OYYI7ikCnU
yQJ8vox1FykomtKPry5NN9WpQK2j+iwyowx9tWCnGtl5zbVP/+k9ryIWUJYLI47U
BM9tC7wITMPV7KSov/ph7CogryZnnGBhhq3YdMf++ytKnJ/Yc6qERixyRhqhMdx1
2Lfe5iFwA+5M9GUNMIlLpIT9JIVT+z5pa6A9iE6d5VZ+Z+g/I6l+D+8q1o4utIBl
FGYoOiaPgJNfB5Gi1rln89flutc85/mrSE/fuyruLoJJVUOvFvBfcmT/ZcANwKjr
VdUDjhTWKBrwAXPmterb9NIvIrRPssy7LYFxMwYkL19LDxrY2T5OpQJCSz0k/VB8
5Ay9mUzedNFoiTWhyGLmu8O/tBGHfYnmr2wW2xS1KGoUNhm3b18CsR47bNLnPvIp
HEBShD/7df0Cq74m0LVsgndIvsSTZ68ddjBVUl4+HNm3nqYnRT5tLIc2JbMVaOmF
AQHVjHMjE+8HhvqK5C9sSJug1aI0F6crosMeqaZiJHOn0O9FxbzY2MzbCyCoJThA
QyIwcWO1azOrJWwr7hZt3QJMc+3DqEY0q/bm6tpDC1NDJi8DB3g9Sik+c+VnRZYE
JxwylyoeAsNOXu7oQXvzLGCRwUlkDr3gvI+BPHe7tbWK5Wg6Wtr3yU23noWPgVIq
eKHIs/eOjlBGv3boZAdbrXCd+kEDUUKhTGm841fzOF+NopEClbGTQQEHK79e/z9Q
gVUI+gMv7IdLzfXEvjqU9O12DtIecn3tGEmoxebGXyAYqcdqjJJ899itBqMxlkWL
IN8A7kjU4ABLGlKgiE1P7cHRT8w6+t3i7+QbiypO8y/XZmHw+R7/nzXYhAFHxhRf
b3cxtWCxCtTToTBAFC/p6XSAdf2Rpfr2M9XQi8nYC/UaoW5mmjWDyIYpRZt8tI9I
ECKrYXq0MkXgVcvK+nGLzcKfsgC1xby245GxW/zHCSF8cpBhlvi0mVYRj/ePPNcF
lYfmsdBl16g3+FKnuWKkOhuf6DfoqotdCpu+9ry/LhTCRiTs40uFHMEvRs57AYAt
JKqxuGY1jMyQ7nxPRuBbmYndAknQIZ2K/CcLrr7nCi2tgjeCdLwR6YuvfLJTEPec
755PO2l5qTfCItube37UIxMV9odJFe4yLlGsikJrIxs4liBaCzbJelpsTUfE3vPW
miBy0ut3pyqzl8yLjfoH966dOFKVldprkEaPWRbISU2BnOQsKh82SWRz1PfsDIrH
9SJZ0pyEm4Or4dbC1pJkkKMGHkoPsOx/hI8SKvhw67qisaaN5Av+Zx1REpGMk3OV
rO0t+J+x/cLkvFlRoSy+n4kaf9ulFgLMRBZNd48FyHR7u9o7X5SAvTRoeQ5RVQoa
YN5Zxzp23jfZ9aIur8LvnSvomRHUT2FCzESlWKtzv5CslKph0NkN22ZJ7z2KoISM
VAUckaO+TbIe0Zc5W8yFZRUm+MlXWYmPCibKFS4en6V9tv3ltBzcHkJjcT+lSHwh
uI164AfRe/YQEyJP4JwnaIxb0jQlk6y+gpmeFcpt+FXsmO0p3WnOab3VrvyMyL6u
OMzuqMjr5A74U3LCQtUDLlN9MPVCjRpLJpxsSbMKsZ1n2afbZMmWe6EMLfO4brJX
gJlj8z6DAjiJVtdLbzFGJU6nl20qK3Gp+Xe1t50oytH76OIERMh0irJEg5C/L3WO
Jwme5RWULSH7y9W+7f4hlh5sll95dqsPXaJHYc0ToXSTJhceCVb7qzTM45Ru9K0R
PnjKzN+82LFfF5vDcIifLUZ2CPkWKv7WrFy0tWGPs2SD2huDmkqBg54tIW4tuTx6
j4pRm+bpveNfhROLnNsHEj4BTdWWPNAzSMX4V3N9EPzlhKizPFn+3XYAzBz7hs4A
Rm8LEVybl1tp4B7HK/O2UARotqaTbb0HXDpvdzseGmhOAGpv9Rn7hm1KKqEqfBqx
+MDnsbOh0CgdEpqmN+AJmnyKRObwh/epxConS1F1nHA4IE1dCJ8IFA+EHAr9dOVo
IKWeljYvRktgZceZXTKdblaGhRPFqdCxaYbYon6jxg6Th0Qw7h4DWhFO8zbv6qxZ
p+/DhsfxqImXfImTIStpUjVsHtYq7KcBgBNJ++N4cDfCfUcaQSUl07nKVcKTsWbG
4M0v0tZLHfOub/K0AnHzFI3SBcwQDnjxElmZCMWFqOzVVlOQFjlcKrfAPJ4lg4RR
OASeE1oewLnCIpYknBrkWwVPLPYVBNxG++rHzTmoKgEhYMQJmw+ga2b0OUl34yw5
ao1J8/AMZVOSChrZdGM0yXF0fjdIyGOogy7T2gwTlJBKq6K9CU80ZpkUTv3YiYRf
rcCniXYMINFJf98jXtOEZbAwLqJUg07TQFNtXo6E0O25QIzWA30Z+uor25D6matb
8lIdpobhqlAM8aVkEm/sWK1tAaJyb1Z7LNFZxYagQGKsnSGgZGCl1a1hqdPpyhgU
6tO/4AfTFqp+J2SAC6Uu52InnoUZYfMZClIyLDAT40MeqWzrWi3GhH2yCgkYRsMW
5Nx96glRy2veYWfWVlwZtenVzx6c65dPt4c+Fga8wkMzchA8RYHl4nTDmWkBu1Gv
qlA+PTZFr8ZiMWLLxL5aP9PoXyNqCAMJ0IILWLQqyQLnkpWTmSLy8lyF0tzI+AMQ
UJ0eCMmaxg2eKVCHcCTgFWSeXknIm9/uC5AMvpkLKWNWPxx4CwMvV13vMeV7y5YP
tsmmRarUy6bJUHhOXu2yjOuQ+TAf6OUuCfWlP/pnGM2rwon7JCyNJ4OCJxnOcYPX
2H/nmZ9ZoazpJ+grj86mCYBzOWhvZrEsipUh3g4q0TY9qtMKB08HbVSbGzDWJl11
EyI0AC1k/MKaeDIE3XT2LRdX/pWudCkUBxwmoKTG5Vck7PyNBF8epDs3J+k6AX7z
IFEt2ED0Qua3cG5zmJG4BfYljmNHtl5BsD6Mp/I5oJzjDfsysM7GI/0PYb3fnXhk
TlGtjcTIjj3Ku7HEzL9B2ihcaIk4U6jH0dSkw0RSVVarnZF36g4TTBAp0GtZjTAJ
dRXXOjDSLFhloXbQdIgiFAJG++a++dS/BRMmQfSSn8f89sQRgHYP68qMY/dhlViH
tbcIJ9H/R4c20uuky87tlBCeyPv/MU6NdmM1eZyMkn8UJv+JNYXfhhOBxOLo79JM
ZLDbA5xa7mTuWAHiFhIqL73SJIZhvVG9s0kx2uknS3AyNOp5Gzd4hph3LHrwTfiF
fl4LN6+3ssT0S9kYIkEZlK3uN+M94m+zDyfQ8NfarL6iVYSQVdi18+meAQnc9MXS
3XbjvXy3q3qiYatgaNs+kXsu/CVvdl/OKDOzrEi5h3GN2zpQbXYuS6oZ4BwoUg82
Y9P9y7VivsyHi+U7Aeu7Cp5lndWoc3k4JKKheiHIcvZajGYK4cOm39KBPWkQjhGI
ijsDLGHxHZH7p1+tCAfr1XlPRogizteO73LUDsNy0rVp/XH3gbl962TovsvfxFCy
qmDCsutM8trrWYsN4gMYb0tqVeDdhI5/aYprDfl17+PdPoyEPiSL6tBb+mv8yVJL
Tz8WcObFij+upMA0P0NG9mdAzf0vZCzigWt3HOcPijb+oWDWEp3BcR9IcOQFpCSW
ZgV7GWG4Q8rtH41OOCX0ooDDKWZjD07Uhf2B6ctpV9XlWm5Qf3vJc/E8ui9RNq5Z
cDxw+IsA2/cbHuMy/GdkZSNpyq32iO5+UHW9XMWw75ecgvxyh4FDXnyZYAUxajx5
B2/d8IeNNlCUEkEfsxVuvQwvzAzajhghv1KZKZxbCO9LnJAiAXkv/G1weh+h4h+T
AggS8LnEALnwsaCpwwh+B55sSsK6/9FrZB2DjjOVbn1zuySVlK3kqyBZPn9fhIMH
/WZP40WMVhzZXpnruWrNd9NfoY14cmKxepp1v0U27hWAGzUPZnZlTTsZZKjC1B8z
8cg8M1RmUlcy64zTvRCX1cAg6rhl5h/eFs6go2RASFnkt0FEObrL2tttC0a1agGH
VUkE9yFRrQ6eInOxXcAhX7znyG6j9KhWUkipQPUvkDgGexjjDTLfmy825KtFsLEM
PI81BuHiwgAe2jGvZ6NBtrIfxy9GE3pFjcaN0se5/er0UY2WVCtgf5YCSb4asR+l
tbDHmCAZ2x+5u/pdi1R2kpYm5PW65uO/WLjLr5R5e0bX2g2VgWN+2reh0Lgc+Tcf
4ZXmdkku9Nt+HqptbxKFihMs+amzB/dYpX6qpFhdTDiuGWWcr0JzO0MiNtbIAdT2
9p4G5qnhlNy+/AkPuTG0jSK3e8jsX32sRy1xnuqd49BpnMRFlnqw4wM7tlS7tx/h
srwfJwfUnWbeaXbz1gd9q4+LQZRGJObGSH12J5ULnwB3wsJszHtVZuZ4zUhTeaxb
jzK1h1aWB8qrWywLqPHIdb6cXZZdB5jNwNHpJPmhzztVtgTqmtxOLgh8woOfLor/
XlD8q1vzsp2FQMMFHJEBR4gGfRXyILNJUmlver4xIf5orx6gjSjZScoH1Bcu4K0N
nhIViWB7tqNe8LqQxMOviUx9bChOQFvAIaYhQ0M1EfcOAgtG0+zBJS+lUGwU/glI
IKYiBGugRJQ76e1In8IMnGetPmhvvDszcRlYS7aVkuMG2ru8lwHRIgzCwilJxj+Y
jhEgCXBTi6p6vuRVAdeL3cG16IJ+CaAdY0gmSonnHxQtHxHvPOhUsPmzobbIoVFx
a2px1tDDzSJZlZtaw7RleQFdTZC+ZIgnZdgfmwXn0/qX5Zw7j5jKUKrE+t8O0m/z
ENNLOnrebHutfyGxk5ztfMPJ5WyrFCmfJQO/w0Jkh5tah7suqhODjUPebZkJxWC0
M77qZEyFH+E5jIjMhVnTy1KfLshfpbgFni8yGTg/IPa40k2ivzKA2ISm7NJvi4Iq
MGh1VpRKv5Qym3AKzjSHSecgKaTqPCAS+zoU4wzpxJ5Jh4F82ix1HUI3iUpEqAgk
Y8NNHnvJfBAifG6CJdKnUl+y7p2J25V+ay0ret0ThoxZxMjMlUY3pwmqyNsCkK8c
tDQri6oBPhL26Wt4iUHSY164lGhOZ1ft8Ewcal3Mo8FextiMEDLHmsdpwHha1Ptz
4zqR6iGubr963FrWc4OEW5DKNwMCTHtiojFhIZKa4+Yee0s5hAsN0DIj1xAW99iy
aTwji8KrLZrUcrsIuEYcDRP7GTtKIPestee7CQVyjCZgEkbBa0jhp97DvmtA1vxy
howYOaLQuF3T3k2ghU+VhxFcTdaRib8gTwXxARzLVy7jnelPK3b55KAdt0AdV5pO
2IeAQ8NYeizRolxMan/hSmnYT2NybZ1rYZ0xnByIISzVctKcd4QINH2lNUDr8nc5
9m8AOjBXcD1mpheMmUnCOa1bPcxkFySK3fDkT3cMr8FJ1qWbYIMJ6LbdfjcT24DZ
5onUU4+lXkv8wd0PY26gvXOfoc441izUBZwItMVfQMfMY4bDhOG9U7vkFknl9Xck
2c69FfC7HmhhMecxWqn3IZ+dd/m2NTO5tXwoT2jw3geiDpT+Whll21QSxfWbRPJU
Y7kSNVtoQRWQ8Pykw44wuSBcpz2J17Fj4W55g/szvzNckCMW4vLCHyMjiCgyz018
UzmLYBKbBTldWdXLGuaGUX9kWR25yMEeGiXL9zQNkmw5drWxP9HbW83tyFazRnCr
XC8N43M20HNuFPHtJU8a3VEvkXso5KppOmKT6dgE+IiZWfPl53lgoCynzafQtNQ+
p3ImdC5EU0t1BbPfi0wueZQrTjBee5oHzOs8LvmIM+90YYRj6woCvaQv40UVI5T0
rMtCM1aJqD+cq22nn2Ax9F7g+HwawPpdS1/I0tUZ8KVa++9Pz2TywdiF4HkTLpF+
KPTl8MOy9H/iTeu0wVxdg7mOiZqGtID5oj+t87qYou47oOsG59TkeNKJp+GURC0N
ZeM183czNJFLbwT057L5Q26cmkRZCCoB7VO4waruWY8MjnUeqGlWPzCMJKxsdbvE
8Fygi37NIgb1zG1kx+VPSaK38EhUaCmzN2HPRQLYyBZZ0nBi0KkvFnRiX9y4GT2x
nxqNXl+9tswI9MQ/M7hFYkwPH2Ei1DgDYc2JF5KCnotKvRMJN/6hbyLGku37yppY
4TVojUjztHTJgGTGF+JcMjkdJh43t22IY7f9mn8PFWoGZT3BiSnwFI0716dZa6rk
OE+/2/bdfnNbDVKiH+RFGJiGi+h/n5GKK3wl+OsvL6e1ibuVhnoeLTXoKLo54p39
ECZYEbW8Ho1E4xp1jtHwFAzJRRh7dzGwhXjuKZAxVRcCsn0svfrB5WVVaBzoY0UI
htxT85Qabzuaoyb0mk2dO08fymmhkdN+uLLniLBrCxoBYGpN4VAbnpL+qVKJom/j
J+QalL8fCLt1DYFVPR2sQn2C+dGWMAQaXZe9iO32mzoZ/yuluG0QBnLAylvS0esK
z/lVMsJyUkvooNOJpVTSuksBcQvfs3pF9i/12G1IOYKPmuFXZMwt2iDpZqD6vtc+
sRea0G34xpyiLUW9bWD5geDp06lYDY2qx/PyyWRIx76HxFvfA6xaHN4fzk3gxb/i
OT/EEOMhS+5fwvoXsF6e6IiVFWDOD9w/gILaXcVPdYnCCLDnGtE81e+ShaG7Xyis
VThaSJjYtnxBpQCHSx7t3LU9uIAC17eqGz9kjOkUf34mwOvi5b+4adbOhqJi2qPH
L/1fX2l2CJZOz9w4K2QANes4+2VTXiCGG/Eq7qMx8YD38taFo6c3CDNLpypL/Hg8
vZ15BpXOVo6J89g2zcRjqYPkxpxO80BfyLnKXm9wBgMfJrqyziVxCM9M1W9M/uJr
nGHxfGlwZJmiw9TS36NCDbK3nTeTCRhT8co+TSvefJd9VOwm60KQyC8fYqsTm8JC
5jjoYtXhwhr7l4SOSujkjxGZzBwuA8ZzeG/cxmBPT8IVyedgHP+ifWy5QDxDcQn2
SkKbM2qesEOE+klZzEfc3rb5Zok3ooXK6llHyhVsoViUU64dW2/iB3bnACc2ascJ
U/GOI4BT/p7MfvYOtGhBTg+ZBekESvIlSRcspRH6s3xnutgsFAyTYh71vy2wWvqN
qHt0loBH0u5QbN5KHFqZA1FZrIF3Z4IcgzN3B9szwOJndXbCZCFezNLB4DeBpi3E
EkuSGTdxlY5JdKggRlbhZAGgwa7kh3R8uvTIWb9tFBq2WiqZ2NPF/JkYX9JjkDtO
WwY/SYzYcUdIabfBLRcaDWTPUP6ftxkyCCntBz2FeHDOIYH4Z7DpKUkm92mxCAEo
V0l/MYh7zhDWlS7ouScQ80i2qhg3Qlk3nlpmu3U1tuGc4rRsqCGIi21rXSXQXuS/
T9OLTfT9GxsdnNds9NpsCktHCF8odcdDwyyElM5QErImn5FFhGGJs9R1RZM4tA0X
/wkQdSiTmTOj2DogojQGvaOuFjdjO08YTLZZEfiYOU5D8/PA0Zu/35q98W+saMYU
UULsuwUa1UtmGQ/4mWMF/NYm9kFca0zpuOG1uYf7WTzf9HKhFerNCFTE99t63+TE
wBeMRFM39Tzk95ASGehh106y6kb5/SkjaSZawVVyNDRmXbZEJsUYG/zBhubZb9IT
KlbUel2ohEYUWid3mNthpXIoWqxEE7eWTwgo90MwirPfAcSh0X5ljJn4Xderr20L
1fdHiHSc9ZkLF8820m7GPhiY+H+YyfQaPgTI4zS7LFOa3YXKXCnM8HWN2tmgwL7G
mSpC7tOXhsLX5rbVj20vgJ3p/vReZ69sZLRJeH4gEorr+QPN8d4qFCIwQvtPkVsE
bAbsw9ELymkxcoeQ3+UukKgERO+KNKAvzRFsSkmyRZgWZKlCir5Fnt1Jg6KJwAb3
J8jhEQ8vXXM1kSHP3ZxEv+dJDLSaYIJ6WwKVUk3Sw4+OyR33v4DFCvpIujlTbzMG
ZWzvANPA//SnVRXqcN3gm9dOkld4Y4EZsdigX89aBCLkLSAaEXX435en10oU6ZRN
RBq9AWOxPt02rSqn//lP3xZnZuhGYOFsUuNdnuYvGxwuQtxijaoUp3ix8ibQM/UK
VUpa17nvJ/fcHty9yzoAuGn7QWoMb4HlgrttXQ6lhh/aTwQQpgQstigknAWi2Mv4
GYsdtnaiVYy1fdSgmq5D3R07ylFzmcNUu+BekZ7rPcIPUP6eWFTBXHiZ4Vm86sT+
bl7IqzWa155SRGRys4YiEOgvoBGMAhDE59f9LfTwTg8RBRVUn44UiW2gHvXBGY4O
GFPuUGmm2AHmH73Q614JczQvRfBe0eyDULhVDAlZPrvyPO0Mugndkm8YkLUa4w1P
IIQn0xe4T5/TwW/8R54oUKc6jYD7rR/jI5DTyEmdU4ZwCkqmhzHTCK8hu6nG/Ud9
pXdIM0QFeqeUTa3h+aOUDk6KLumseYq7nt/fcOWgkuf0XRTf3G2+R9nmmi30tIX7
e+xRErY6I43ZIp9UJfCEyGb5JBFELppXXUPexT04j+P+Cw91oAIhkSzQQI93eOx6
NM8txU5nh5yR6Y/4J0Hl7nypR1EqpSBIikLMGeLfQsZhujPul2Q11FPmTcBkO64/
CP2EbFT/3g1LeYix3S17RlvFOx8wmLENi+X6K0kA/K938IarR6dAgqpGFlxjw/nf
viAKpkacgVvFMz/TqtTtVCS8a6Agx4fWJwcjr08VPlYG11FHE0IiuDChy1ZpNIVn
hBbVQ3eTE1QxuKrfaARzx8OH1xPGJDlN1QqznTEuyxF1ceuGc64lbnSD5xVJ8NFU
Y03b2YGSgOLDUYdKFyM5YI78RUP5GRJTETvcwXvyj0znLI+ulT0bct3ILKPnBz4h
A6iGMXUqZYc8eG5uu4GcrNE6SyPX9xAjCifQZuCy+uFwRf43HRH5lEnhv4y0efUV
Ze8Cy9bdv+DST450fvs0mOfII7rOXahzSpNm6qAr9Z51FmZvfhrTT4jq6cgPAE37
LO9eVHwf+y3SxW1mTRY3REfUVomDiB/NOiOdU3dXXnmgrnW9jZpQ8T1Oh9PfgAxc
O5D8Btr0Y9PzeNSb8NePhmK/Yk3VpIrnG5/UUybumIDG8QlLXqU9pVvjG6nCsuK0
ecxdYf1AI7MFVxMdFcZ7Nc6L8Eipm0UNeNR7JwgZs10+kIAEqMUDIyiIDob2/ncH
q5MrXlNUiCY5qaSr2u+7cjRr+1uKsBUfAWZvmgRCRhKN0LSJh7+y2NJgwgqkd8ai
gUylmhLjMG9scGOIjddriUGSyZTdRcYF6bB6UzN1E1e2GVwKZi/dyKs01WrKu8o6
aWKufTmMjzylNuRCGwuX7wMkpFy27CWQUUqm2jtROCRudGVIhvpqgGhKe7xKwLhb
bbCB997pZXMUhhO6Wh2TEDbAg1q3gJzuJgGUdwT8KZ+rWNc+MlBQCnakf9UxKWvO
heMvaYzJTGeQw4ZPhyfuK/r+k6TfJv4zyM7Sv2T4PN+BuPo0ZbuGw5jT2ACZQGzv
IOiowGJseV/HgE4nTMEL3itOcBjhrmIO1Bdl1/0GD996cfCxyw80Ia/MwB8a/31J
s/3352uHryVm7b2+OSEQboHKN7efRFosccWFS6pyLkTiiiAjKInIW5/rap9p2Sgl
RlFM9gDtwgYYYv/TXzBiCnWKjbUH9dOGdlPLcAGngzmPFA+x7iQ1IVO/yVcmL2oU
54OQEq5zg6x5rZem6TQ3smjvjg+LHJhwIGLl0JNoo5Ft3Gs+BhLTxEJhR9oP4Uc0
V5hY6ESVg8L2wgkd81F6jmvRG2IXomOrJdoMQcB5oXI4Xe9i4clH+k97eqZO/OGL
xv4ycsX4TwkxedbZA0jiSLx8QLzMrIUVHkHERwzwyzx2SKw34oazYI3P+44YTjCg
s8INQTp4CgTv9PYIavK3UuV8HlsfGUXOcVcs72WwGtFUYnzeMjwws8KV9CGlQQzE
QPFXVDpgDP1RxrRLiNH0Y+QsjjsFhU1kBd7zkDC62fh4DwMmSdEWcClMFzxz/1Qt
K1UJEO8wcH7DNMsFQaJKmlLlnv+Q1XKGbgh6PQTw2CroESy8FYHgDBmOmNgpBSz0
HoPf3QwgR/gFylqK3jTNQkJm4U9UEpK5irnbQ7ktV2xTYs2RP0upcNeW+eeJM/fx
vWb+QeFMuzAyw44faTgZsZOWOlqAPAYgq7nVFVVCEjq1jsIi6z/QVoClEU6gwg7i
MH3W2ORdLRfELQJWKGuThICjfxaKJVBs1RS+yb0iVbbT9SsY4e7NEMuyzLyBSIXc
tk/ZbRinogaty3rhk2flMYK92XSnaZE48n3gOo3ZpyMIpHQelpDecFnGylwDg6Tk
CvMC0asJDhB/it2sRfRnSxYcGmw3fyMUVMAgwFDK7LOSXB9VZyESQ0F79JCrRXs/
aUpkCuW5MvTDV/7Gi7ssxGGww+J82535ads9CgpbxWSQOQKGoLhj1+zeWC07JYRa
bkMLA86IFIwdsVKjoZpObDkBvOqExSMHvGWGtNAkd2sQMH2xR6/+2kxfcO+DcZ9e
rQ4jQPTjoS2CPOdFxN5E+aqe9Z5Oi1bbXw/O6dSW0yl22lCY29EF31LRrp1pLlA4
m7F1kSdFHIlMY5W4pEzxVos5ehJhxI0dzCeFL89N/nGV4uqGonKNueqKgunNL7kM
QGdHoK4Fvq53+aHa0zKexe16XESHts3vnzJOL+Boo+iI+D/iUc0QJHStWAk+Os/X
59SHjKNXfLAsa3JuwrM46qCRvsxLXZCm61M4o8ZClT4Y15beecOs3Qd0NSeHctfV
UMwh9Tod6HXM8v55EpbQN6ik7+as0y6j+fbrF0dKeN4urHBJestNDAxzny7lBrpe
3F+surJtg08n5ZsjAdnj/tte392lme47BwiLEyd7jjCuaEy14+PtjL3iftJwnywr
3zvbJgTxRy9AHl14zG2Wp9tjOEtAIZZXHo6DJsK/p66zVszY6Xm9jvIXFixdr5Ai
61U7AG0463H1Stt6O8e3LeMGZsNeLJfUrOJEhlSEN5uTQuThBvVJs2XoJIQ88ymW
gesKrNDM2AGwaE3mREJc9KuMDgtXlXOZz/thMvU4HtON3tIjRDO5Q09ZcM6LfehA
jnckLid/K0KtkeQDXwPnYbn20zZkMOtTq6TG8J+AJABfREuo0ezfCL1iiKZ9XxxM
2EKnUE15MMNsyF5ijjspG7TZjfLIZavM6A6dYzvA2Dp0zip+CVRigMy81IbRXVAp
d1d9sdkED3KOv4Q0Q+srO6FrvxtE4aLza6N08zfyQc2Pw9y+stIevr712QCcGrqL
+j3W5leTASJlFUB10Prt0T18nRQ0unl6dwLXIjz9fp/KD5756YkkRTPnhjQ07dFA
1xR4QKCWFLpKP6gbgnkVJ5kjEv7EJHKKamxOGjTXGMpV5PtRBBzF/xCi033pTm/0
b+e31rEBV5lNs7OWeoolf7JIhRSvPu+WUSIsDGMXOs6WQIdtDipFGeP1fB1TjlRw
kBamI4xRyYthzgtHgW7RBRuEVRIdkHfZgYxcJAXqRqDeNB/O6Ks31BNWtZC6wJYk
9lo10/m6xQx+uRtkbgPlWrO0jGS7Q0RNJqxRYwDTyuCJ05eAd0ULNib4gw/nn2lh
dbqYZZp1q2KS+ySKKP1Ox4A12NfCKHsCVkeY8sfNoVNciVe53sg4ndpA1orLCn9R
wGlcp/kAWX51Dc0SKMfMHMWPxPECxm/iFugudqbS7oZ1S95rXxNGQzp9ZPdFIl/Z
09yrE3DgSfuWZGBGUbh9Bpt0MwLp62BmJC0KBLvfZW3nsk9dzg1Sw2ecWmDnJS9a
l1fe3cuXtbpp2kStxeFpxQZJYu31ITOqhRgJ7HPoqcMZJQrXdZldnBWfW722CoSd
stNV2wW3GCQxXNeRIn0cypAYN3vPrPgPSJnj5RYvluJBNNpjuv7KuKDkVMiELeAZ
+fRGBcQZn7fCDerRHR/Kcohc1osH0Zlid3u+LnnFoFvfFdKdBILxQAIGSoC5u6iS
2Iwyp9NEg5Exr/VFN3sUrWuFGQwscfp+Aasf+9VlFw462EMkbrH4aG7P5P/HOsbg
9xvr7EY6dVz7cwJOIR9QvYdk/vwnNiV7FoJqZv4JuUAL24BZ+y/9Wi0X5hUwpHEQ
mtAPYoBSj+Yg/eDPNuNoZijWsJoyJcEKNWfiCpjQSCmBVOMHZOxpJoaukMmbiehK
a2dnHWjvRvO5tJU0NGNZD4YEW6BmHU1fTt3IPbK4D1/Zqhjlju+OMMBfufxrtn1P
ph70f8QaBfn2ucnMI+ZYIadrkcFb39dkhLmOvLza0KZ4a7aN2VnJr76EHAwuc4tL
a6LdmQ48/+4qsQFbiPBEXMo5A+P59+YYJ+al0yL3hmFcb+iZgFttEu50lV3R7Wt4
zyvLrTMapr+1Ff6pQs6/On4Iuo1zGEqRxLKUQhhMYsTCCoCegKwJU+kMRBEPjKf8
ZdvR+24RZ4xRX5306VLHTESAD/2tULRBcyqPwi2W0Jje84NReCOell7eSedSmp0x
RzzkQvP5uhQYvd2tB4t0dzb/MtCZ2iA4cL28+tqD06M7m8XQMjuh5dyUXp4c/rsS
TRTHpdPWdliVx0XwvbEBXZ1zOTmS8eqJOT7AoDffkUeibyQENoS9sdOXNU7O0MfR
qwu6x76cKW2bGi/599SHY3JI6EY6UzQQNhEgWLcUr49+40rbwDZNPNTrCd+a0x0I
+KyuHNe/2WslmC0D/pri5JjIUkmp4WqvR2Tu6QJevS+sOk/2nolR0D2TFmYlMG3C
jztKlxgrY2bLG2Gaiyo5sveEF1LtUK5T2uQO2/+jNGlB/Yif+UGBUW+DIZsoOXEn
/ilVboGRHkU2QLmTvhs0KFL2IJ4uy8ams/fTVFGUqVi3NWAM8FprrBjfiGtaUq8h
d6z2+3KINitwEpZd/BJDef4PdtmeOhup8gpzuY1Y4KchQuyFeuINCakDugr96/ZB
6Q9nLt8BAQKOvtTtrWKSPFNJcgJP0l+j94fpOw9xmXGIr+QYvTG0H+3o8i6zNuRy
i/VYUDeadsCw55U/PVHmEmuavGdUZNU7uQu5Quqn8gaMylDuR+/ZC64VZPRyJGEW
zIT6skoOhg6fMLJWrFJS5EFMoExw1SJ05cnHrCBnwN5iwqMVGLf0FUaPdAUK+Q4n
NkbXbaLFijAi6r2RkwacItmP2vMFwvq1BXtQyF3978paofBZObrWaoiqsxnoTZvr
ifRKZEPJUTWqkx+3ZgAtYkKI2tES8qJhxs6JIDpN/qTLm0QryFtRZMkhp4IWz3PV
3pJFpXhSgE/1TeqUnWFGpGek2eyeiwp+aQhD6BpazFRKFccQ+RfVKWI7WBiDLtIj
fsi1EPKNn/3hmJj8uYQk6RdSJLFTACTn5Mmr1TCCEJH/Fn+2FlPHyKg2K0BFDXAc
HvkLEAtqxrgiNGGGizRHSkektV8FWhhGiV4vKqlccdfNqDh9UrDqPqAFvqxWUunx
6EuEcElGelDMdY0jfcFrtfzp9dJdsc6tR4blFUKFWyZOLgLsN9stcYl/aLJetuBw
1Osiyde7MXNyGE/aatXUz53LqXhCv8/h0D221XHZRvHeFj4d5VDl7nn9oPPzziqy
OrknaUsUwsxBLgGAsc7tEMNLTZvR9iLXpOt2Yy00MMC1lHNdcbADsSKveY3G3Knk
wd0QIFB47/KYfRXc1qKHAhWmH6Q0K5golI6rMDz4bEYdq3+rWJkQ4o379haHALdX
OaNjjfCowI5n+PKTmaQ+behtbVMw22X5y5Z2L/YE0spQShiid/1YTG70FAY8lPKF
vVHvG6ez4IVOyV4OwVtpD1hJvz6xAIrK+hWZcpNRKgIoIlyPqPYPDjUoclLVzEQb
k2mYrBxkBqJ6eipXXuMuxk/2HCb4O/Ql6KOo/tWv+vrG5NXOBoOJ7D7uSWBEHpql
BxXD6Xvesz2GiRAFS7yfLC+LFxMHzGCX37yWRt/l+5qZnI56+OyI/2/ffhtddVTJ
3xD5YGs8KBCoZOlPJHRmUoksiSlcWaN8fLKK1RaXHTZSwvBuBrjiapxX22xhOxyH
wkD29fwMzIrtVGPkLTEWOOt3kmtJzj+W7suKgkXhRLgymSyra4zvwSz8D5lzKH3w
1SqEi8i/kDJNj6H9S6cGWQ9dDOGaTK/NQw+Mw9iJaSYoEVk5XBCvjmbWlxliIeoX
yrAypICsLCx9fs6fvNkfAUG4Ig2s923T0aagdiZ7ZlzC76InuyyGdLbs64CBsTU4
Fp825El7a3q7R+c6b/TrC4lF+M4YZCPha5lv0NckIL2cEb8Y+dFCB5uvti19NIdI
sxrrfN+qOT44+uxYL0qR8mwy60L9314UfK+P0c/36v2Cs1TxrlKMPtJ98QKUmg5E
XgxeDLc4YDNb0hkSw6dr1jLLVpvtlhestEnoP05CqqrhdBlePFNmWXqjl0CSIdsi
557dwTDtVkjpfW7qn9c5PpKpo+i/KgncfApKwIlLUOhpzpyVocpWtvla3pYtT123
sWCt1ghiS2Imn6QIFZwaY7lEV9/9XnnUntsi5O3hVmehRKYU7tMs5vKNYKCCpiKZ
dLnp4rGK247Bo0vagKBVqRU64Yg83VZOtILJTZ1cRf5rCdGJcG7a5SssMGZIVqXs
3DCRgx47dCUSFIhgPdm+y7jPU38jk2SNIk+5HMIV60N463c8D4GCdX5kk+u5wt4V
76Vg565FsLj8m+AzXz5eY+a8BGE46fKUB5yczRhblaQliqUN32eSuSBcf8ZeKiCn
VOnqJdfRpCe5QK9s9jVKK4TOQ4zYOO7d67Fg/hHPxPuT1HSXpDKRGyU6J1miCiED
jP2AnjKyxRBpMIh1lAXxJdagLsL68r+oo+HgoHCUYBQZG6SkUNDmN0rQTxKOGUv3
wp0NVukpoGYsrr7fudWCumoDMwBBUmoaTxqFVbisPzhfKylU8zWZfn6iEOOdxMI+
VFcWNP7W9F7aNljdlwlNw3HotZcOc1t62TX69xLEHZV8XSo2T2q/i+DpuWDf8LU4
sBE6WG47VgGsj0CgjncuptY8tp2hcdC047gJlcK6aFnLDvLSqoeu7/toEttWfNFl
OZQcVFD2eCijSLuQtodptwW5h9U/tpIU2ZH74SmnztVZ65ucmksZExnjzA6c2fnR
2dLMV/69z95b/GQ3Y7heJjPLHhEDU8ZUYSb6AZslbzx8Yy0OpaQ/nd3jz0EFPsr7
leZX9GWSK7TyfUFlhBb80/5cuE4taTDJn5YRsN1BmlKXFIrM4onVPOJH73+6OTfL
CZ2Rm51KpcnwLPjJeP54w2W64ESj4x9FQL7SlAVpYb9L3DFR5tNdJaz840oS7NRV
Sql8APTyRyFWFLdmgazjW+Dv4fS63eYFg9t+TDOlrZPMoKJj2qOaYLjr397jDQr8
PAFGhc52d05jS+cJ4UE7kUD2p3RViOohceKfNMRFLM4Auzr9AiZumsoX2A2dEHKZ
4geyrn6GWX2Jcic1ibi8ptyPeVjHIPWkTRmEdmaAGqaxAudME2ctQyF89Uqk6Ptn
Ot/rpnvWXqj+YaGq2RgqNPboMFUeI8uKoq9pM35G4SxyM9kgxtMKGknBrf5m6N6c
HEQ1MEWGW0pzppzpdFfrRyZMPHXu5/zsWxJdLR3qNj8Jy3EilseZOgyN1J/bXdHd
X1PwATFG8b2oEpS+qEHEHUSB1pMycO7VsgQ7iuFWYZLTNUZxNLMpgief8aYIaI5k
YWPSDkGSH/PcF4gglVo2w4vupB2eCPD2ZKd4e0J7kDSupoQyRlo5qc6EMFqlCibc
ibT2V2cUGOOkk6pCbVoEqpN7MmO7NIo0iUK7J4CgwhCDbl4iEgWAy4VPqHCJlKM+
vdvxBUMbz9C5UkztVaOTypcHe1+NuYIwJvmJXX/mHZNYhZBSBQm84/I8bdLYNCC0
Kz86rw63fWUkYOotl5kIYug88GbgKAPSLiK0IDEoOQfH7+OaM6etCguFOrAnCGGG
MBsV0fJGNrRqJD1DOzlwsk5R1MedAAt/rUSwp/5U2gpM4d6CJ56CkibBGux0HqK8
DBZozzLSLO5iNuU27xliczE/bgrrEhrUE89fH9CQmha/7MUhhr8YjimZQQ6Vsbie
5uBXlm8rMb7v5rFRkusBJrWPGnlYkgBbwLbVgwJz51D6j6WdPbCSHzB5RXU0uJ1v
URhilmU8xYlminu9Kr96qXuzH3epyJAicmVE8xNq/p1y/ikQt1H6QICtDI79ool/
vn6Gof15Ugh6JfLqLVg87Jg0H/Dm+3Wi+1omoauPaBNvPZe0d76IcefgAUzBNQLz
NwlkGVvQxDLMuW6Hl4sN/lEyGpFjadkrEZwpFdJkEXDHZe5X7ktMRLJNzlDGbu3N
5mxQUNllqTl8cfB2ZzzG1dG+136albCJjif/DOtC9AmtzInZpqpkp9ATnVAc9GL+
3d8dZw6HXhPtpoZWfX+KBxZF9SGdubWXN3R1uAw2foxJ1A+yKTdxuTkEXu+cR0a5
kp+Tb5XmbhtoevsnBjiz1AapD1LTRED2r77ImIPy4xsMh3Z/P3B5Ep9e1ns784CT
sWJc2+s2CRW4hCu4CQQBLCYIyWWibKEYVdvPGsS5R95kLygX0dTFMEKepjc3d6hB
c31++fZyvt6SMcHqv5YsdnOMo8emUEYgN1Ty5SkD79ynkOIx4oMTiWIKTq02Wpxd
ctUIaO2h+r9paDeX9a8wqqg6zCfhQsQv1cX42BYiLpYkKgfViZLYkR9T7ZuL9f0C
vtVfNYWHX3FV1BnsMPSqwJAQUSe7W475TV9rqQxyVUTB/ThF/lHFyX5AaTP2qWuF
z9vhzjmGC6Vv3ARC7E911lyghsLMKEqCUrlKaLhPJc7BhQk8j7R6AJ8ei+ajkjnM
4HNf8gIyU38VRboa09IC4i15DxAl/r+nSg68r+cEXeWJXbrAFPlpkMIsZwR3rrq1
xvvSQGo9MczxV4JbFAbr3DnIA83ZTQ+QUQNbSTKvB3InMxr4+DrBHNY1eqScrejd
l8TwBGwhfjibp4njRzz2GInHL/x8OL22sjzbUWgpYDuKPVzl3jsFqFtW3kztd8+o
O5VzhsgRLNmn7/Yp5BU0gVEjfTmgWJHaBeiBh2NFiettFkaqR8OzCk7ZvU6qHsRD
PCrzqLhe1UGsx2AcQEIODukKZ+6rcusdW8vmWKkwriay3cfwjYcdAQMIPk4cSCvA
1gXMYmj2TXxJ81Ro5YMqK2Om/bMGsRzwHPr8i6a1JAS0ppZB6LfWo+DzGfSpdpBX
dHEApz/D/KT8GEwFq/HO3zZyCevYf39ZypU4ypcpNumJtwABE6eCxuDSqj8edsjD
pf/Xy0EfAOlOdb8AZnTAGhP+79it2wJJqUDsvjJkE+6zw+Bmwig71rJdarXs17np
oAVJ+j3DX+k5lXY+mCzkkjmsN/Uv48ssdgoho4anhqsnTJYIquvqWTx+FpRTJ7XI
TpmKnoloishFcjvIFbUjN2pSefXJkKWHKAoYoXka5nbeFYogoHOewfuu0pSwNLge
SMLZ9Gf4EJdz3KaL66LjI2W4kee9aHokdnrINZFFiHUC0IYN1t/wW6+aUOeLWZkE
TFlKjAqX+693YluBt/1p6fMtkXgjJllUYmHqbi96cJh60rrDPnrJA4LBN1Cwu93Q
5hlXSdQ8YVzEADJ0RTZuCPev7R5O4bp14NL6UsFiK0FV1Z00AiNQsI5TpEwGvvM+
Pxjsii1XUsl4HfSp0FZfxKeI5mshYCH4U/MuI5we0dVeKtUj7ll+Ko3Kq6jmlDM+
sW63DLL9/NPtEKCRySDBCePD02p/zbtN8hiYGOqQF+gtBK7Wrc5DBuSSqGVRN+8X
hWzhsvlb1iAdOwPJEBpTI2dXQB66KpdlC4yO0np08v4sOsvZRomrAAoTTGnNwGg+
8oagX5oOKyn42vGaX1bi3OwLxn9He6jXLb8STRAlpZNiuMY0fEnB8fl/Y+P+JcQG
4fUTPrbepj06Q0yBXq+KW8VWtqWQEMIxGA9azS98VijWyAywZLmcjUqPsWe3zVgj
H+bb14LbVcsL1Pg9fWQVl3CySzqCbvr3Zy7Lk/yrWs9aQJHsw2rLFB8hwnvXqLs0
6wATAuU25rEtQSldcnQBwgx81+DzcWdGlLwLQhQ1sXP7a8UN11hAP+IXwkHfCc9f
6Ds1mdGPuKFTE4Rmj4Q3u1JfMMEOTROO57kgk0ORwRsNpVGTgNQ8TspJhuA5dqtv
S3YaBwLmMil/Qumv+nbmQrzaW+kPP6jBdzDb5WD58Wmb1aYQhuxL3K27bFN58HJ4
VEDoJiUdXakLDzuCgP3LyAfX7oC3xZUzXmVbuT3mSYyUgWlkooT/+HErXC0ww/UH
PxzpvxVLq+uAvCrM2gccvRu/O0yB+cktrWRDvLvAR9E9gTtiT/D+axTlYMQO3wiC
g1wltxqgGQaLEgoiCUdnSjtirq/bInXXtcWHr/bj9ZtBuFfuKn7AdLGTmS1ZQMUa
4RqNMxOEQ6IIwjEFzqZ0nIYaTq6gAj51HqmzKmwLq4V5I8v1AJSMtnhG9r1wv0yI
v8NIj/EGxgq0soEyQRm5Lk3VEG5PsIeBvV5E/D0HGgs6ko5/uFbejpU7EMbTRvQi
XlEFxShd0+IPlHUAgxfA+AfYULLK/WzNqpJdvkyEbdZUbBw0PGCf9Ysu9IsIXFKT
p0UlmRguwcNpm7pTgZIX9smy+ziFIeNFyU2P4z43L9ATcxp9CQuf/wXNzzmMz4AW
02lqMPazVn1ftxz2wTRGvgYEZwgE7foIZ0ahptRl7lFwGRdQcRRuPY+Ayx9hOWWY
cEDCUi4sLBitjEcKQD/HLA0nu/ls/rpjaqPQtmuw8X2AD7NegQa6Mnt7xnTpo5E4
2K4xoga2PdVLwski2G64CvbTvGFacswObqECVWCz0aLYokwYpsKuvUDse88P8Kyy
VKBfPvp7U7SxPfjAsAtdRpUlledomsUJ2knPgeOAQ2TkYiLcbPYrzB469KnEuqCC
bjKBJ9YKFQAqEtfdQxoBV9kNiOERckDXKIAwx16+pXW4kF5eVdT5Ox49DNmzpNcE
/GQzYrjYgwKs0b0adY8ICqt7YGAhjFxj/T6Gh0Hjp0g5w/wa4et2RHU03iJ1N55+
n8XQTQBHUnsMRs/gp5hIz/kSsCyMV9FU0RuPa68pT6GakRNFuA68r5xvkxdmu0gf
yNyt5TsfkMr38PKtcrPFevjHu9QfiZ/wLAN/8xJ/ZnuSbkn7OXCNHc5CYTVG8wU/
LPXhjR+ovFD3qwi+T6ffTnQKFvDHjeC0oDpO9e8zTuEmzT1xU1V4UekWOTKo+LEp
drbcoPSMIwbSb/LD0KHagfbzngASxE8dxjc2uTYamI9pghKyyzReETu15ZwhsIzN
BMB3/YO2li6KnnweYeiWO5aikiRZhR3lTC5ZwGpduavrbD10dApAgumhUSOri+Ik
Z33ogdV25pFofEnQ2S+3qkKLJZ6MTuXYPpK5omyAdOLsZEvcRsxzyBheuigumJ5Q
f9dhW+osmN9de/W2386i12ktVnS/0u/+K/5U+P7l9m9NaXS9QoC/q8BVbA1A2+Z4
Dai7iuuit9J77by8scFxdoGXuAW5C39WpG5rIvfDYZ+Vqi8xJnWqbcw4i7V2rLrb
sKa12+t/j4ZpvDtUu1SxAolXja2OZuel2r+jrjhTEDa0ASo28Rs1ZYfdRfcV7CcG
b2qj2rLP/M2V/+tTGfxqM/YPJAdtW2ULQ3UdCfouqH2cOLWMfcbCPDBHsrcqk9VZ
XB4BfyKdtTDWynvJrMOGeoTKko8A/a5V7TwKHagDRY0Q5PKiRlHul9PlTHHk9tqK
fguCLDN+g0kt+QpF8vVp86JnlO92MMMMabyLFuhY2XfUoPW2PXWAxWONmZsGSfHt
NkAFOMfT/u0vhP+UYpmYUXSrC4M0V6gGdE36rPJfMw7lXqKNJQ/ZZASHPyM3S/OL
jXeR9Dt/WIvebovf5eNV2N/iP9az+Yy3HJL6hMshB8FGv8U8k49/M6xvFIqRand0
1hp7aBgTR2+gnicau802ewClhv+XwUQdAwHXTsqaoqOstPxwg5Ajks6RPPjQPIwl
48Tb3cm7vdAl9jNgwjKw5u4/VXfyX5PRHID/cgBN1kTXAJyWYJZkLOfQMynvqYXr
eVaQU4l35Sj9Ej3SS49xLyHvK3CrjNmGbcPLb8RIgFId2/YpVgD9uRe8FCSKRFra
Yf6OvZ49cIxx5YIwh0tahFkDiXAOu0SY+ubVImSQN96Xsh+/PvrSskNgWedEaR3a
6ScQCm6c9FA9KGA4+zS3iZXxv5/CarILAFk/g4XDEJqQxoPwPzOvipeJ0mHieKq2
S2RjQFPDqyTsDgzHiDfV5qpEoRvDpBhY/4ELGVuvf6zk9tUedaKB2gLgYp5t4ZlG
afMvPZWLBR9QkQZMQKteGPBS4xO/QZh1tUn0yQX/8HFjhVd9Pj/+/YpSeqmz5Aew
cAT4Vhi8dYy+Fajl6/GRE8zj6f7XaPNinpp7GRpwEAnTm/0FnrlaZCuFBj5lf1Og
Phz8+CmJ8BGdtxHj6AUW85MsZnSqT1fEr5wbPce1N374lNYLkKDvrkI17u1nuZRN
UEM7Q5e7v1dDLjcost+CQRXadws/ni7uOx90Bbnh9v0eIJZ0Nkf2CI+uztrIyCAZ
BSoUJ+yuRFOxBhBnGVwxZptiRtzkEmNyb0+vUU5Dep97zvbmisLcErZaRJnfxT0B
SCzH/g4dT9JJv8dWY/cRTXF/MyKz6k+nFAfTJSdf5EnMU7Ka/wJkpOiMrFrE4wZo
midxSzlX1qhWz2Ty5gg5/evDcsgyvcd12XrijbgMANDumVS6rxOU/qKL2NKRCdqp
GF9CPiEG7TqOtTtG2CHWXc1Aau3hGKQEzO+4d9HZ53pAFhYUZnFpC3zl0QY5CKbW
A310QbcGdBnkeGBkpElH7i01AVe+iyLUGDnaLeM1rc8E2RQZnfMdFhVFJhWvm2py
4evdAdxiMTFohx+JtAcdnP7oeo9qPp2Y6rdffuWD8ccJJHzRI6johAdxTyM/i/HW
kGwEpX82DvaLvcWnByFrhbxynyq/n0oWUd10YJUSt+YQypNwWxzquJGAJEGeKRD6
e8NM8nj4zsKikCHHo+hnS79d4gQubDzDOHQ8mmMJ+3z/dPEuH7fOZEmVT1hQRiga
Rf7xkuaDied/sA9K+NNpZx1mtKRggvaoagjtC5yIP0O5uwlUoBXeD6ttn9ccDApR
+9W0M+3Fg6avIXIquzC8tM4arMb+sV3/CzDMUISAG+JeUM9KRHUtKlHDuFkhPzH9
PgGHNUQxDubYwzL9pBoq20hXdNadkLGauzbQlnpT5xX+uRp8aSk4Kc6BHWMA2kco
ezL3lPNZiA55xjJqZMKdsszsWZNeistvV2oXHofVGDx479Zdg6EzfqI8N3YBP0iN
paegJ80Zp45zfhaFyuxj0G4uwUH7idSZDkudJKtpWBMRyyfGf+FUwkpY0d5YoPS+
66QXhp3U/aaGfedCZrYGMXfdVMQzrolEXBwmHbzwWPSpnRv80u8zUdhjrbs45FrF
GeClzTFOUevMzDCHKHlJuqrRYJdGOmSQYbgQTKP1OfyNjP97WRknHlnUWCj3NZPu
nKENlqFP1TpdtPklAOtGg60cFxwPDmut8MGZLv/j4WmVzaZsTk8n5PqhakuQnK1C
OB7VpEkkOjHi5uQiuORd6fFIuQdMfzG19xB/en3Oed5rnTukKP+8r3+Zsy0kDrnv
HSnLZx1KTD2uYkj4unXNBCjE4KfmrCArwKE2wF8gadpaG+SnYx2QwBdh4l3qeTKb
BgfzW5G+3A23TxGgGWUNABtQaBwRkXilTlfqLb1HZ3AThAWOv5U8yE45Miw4b6ZB
yBaUQVGYUdo+cc2akTk0ucWyjPB+DA7MOi6jxwvgq2gYKsPTas7YNMB4oDxWqDCm
ZIDVnnysyWpkGBbHVcXskGejE4WWe3rjGbzF1M2efzKfbHwTq9cb5uo9zyEoC4et
+nMsh6dKw/NJxcMrgTU4vWD3cQPmMiXVw0Uk4luR3JsAGpAtsmVxmiGacqE0CPch
/rQ0K3OWEIQ/Y4vZSPDYhtwCY4zJpsADMO8ffTOvT0DMqwzpElOAlL3nqAQbsOXS
icJ6iag90feGrCji6rPZ+gIFzaCcjUZZYXYVY7mXyTXVs4iinwDHX3Len99NjW7/
v1t9DmLUgOptnf32Ep0TJdIPKuykH9I96jAnKOPQQJHqt6rKVRKfN/4TzCmEfSpn
SVJ6r8JA6mBIatEQ8lZrPfIzoun78E/xJmrCGHt5bnJHV1hsube7iUkYoWhRJ7B2
kqEerKHalSHZd068PpP4tEtWIcC6pfAmvkhytbz/ZfrsrVF5EJCHeZ94qBhYlKKU
b2S+hyJSfGCqvNmRSxrKONzMT13Wl0sWNpZI/Ik5DUcje7GLrAB9x8Jvlu7cVb1v
AwGbO9Un3Cf596oGqunZtKW+ZtrygjXmiby1R/LTwrYRCDO2jLjxyosQJ96Nou5T
gwlMtzxpGPu6BAEfww5GCFY2dk5uoI+RfqHvZFPNXPYVzOdvSzDv7d12Q+4lyEBt
jwnWoe2rpQs47EA/zVxg3ay8bK01m+xV0t2/wM46GQC4RzYKpqX6aT6SHq+TGjsn
1SOD7gechwqNKDDtlTEDU032jb3cxDf4MQMiR1ouLdxjkEPrq/qNUUZDBcrp0OVg
Kf0uxQLxnlZrHkHOvYP9TDJGlGZFeV8312SDHn9J06C2+OSOy91LgHMLHHZ2x3Mm
oDlfxdSOsnojnNc/DLEWs5/PqcShqOgNyGEUkmkKs0o6mTi0WjHOvUsUGS3LrNSb
/YekW27DWjwFQop4rm5X8u3Lpqw03w6CEyePeYxqU7/ur5ROFoiH+1r4r5/5Iq+s
pRuUKGSWeXzuX12aY+L1PFlBEwsAD49gPzgfhhybX0X8FK9EWt/0gu0Ay7XzhiI9
DdCtv3VjuUnI+CT31jp/4hQ+21FkYdaUWW+5Z9w4xVie9Tf0Uz5eEGZPtjXQm2cb
tr9RHEtbYN+jKADIlM3wmlktc89/ERP6LlxprIOBu3IY4W8e11iE+K52pmACGkjG
fzXJo9R7YiA7gR3UJiYmZSj7IPzhdtA+uiv9KMGlu299XWvdE7bM/ieAuNNdm6Nr
xwDZyzakhXigbQzduIhcxLYTngXub+dzoEIkRuKntMXDE81/IBNXO7sgAHLRYp+6
Y/DLHPTP3o7KnBXwtCdRApv3hDhD7NY1IWYCSrXpcqaOwmF/t9DDq7TCK4Cf0P+J
uvukPnoSedg81prEa9ONOfv8M546qJYqtyLl7wOPnR0J8TAKLFKPdTd0T2FhjBD5
FSx7Oki+Bl+hL20l8G6sjmUNGDln93SfkJYSy4lX2NhrW9S67vDgqd4yaiaOz0Ne
ystuphGjm4Fxa/8azMfZDOLUkpj5Bn966KjQL0pwgVJCXbJz42o5dECRp4AieDqN
gj/XiS5EWbq6Ej6C/XQE4oQpHGSvn7hdLFkosA6LgEEJYWOVyouX4ZB5eX4QLpJa
MM44YdU5TlnX0unp585ktb6X1RJBN4zl515qWImmsyAiVlEntbGUXCr9i88jQG6K
TQ9OaeARxZoFWRDXMjpRzkl83k51n85/v/INdr3cG3l6xizaAS8L0LAuQ9oOZ+xI
C4LrF5RKjBxsjo35v74Decx0Y1kffF6VBzjk49CvcBI05ViM1wLOnO0WpQz027/e
6Re4GXc8/p9jcfLTppvvx7FfoRzdpWc1FfNgQ7coGq54xPO/nompiBPDxDbWq6+W
m4oPdMKPtBEvz5Ej/f02g3rgtzrsk0oDjBVzK17yFvquLSBZHVSWYIf0cG1ypcza
VFtvyIiH6Pt+zbVxtn5SKmmFE9WGT5DSkBzUf4fuHmpTlX6AwYRp6RKCvITtLDRm
7J4N1l1P5mg2NnSMliCZkdCedr2LyrnbN5wwJuVlzd9YCPjTaJ6deXF6V3CqTmrb
0mLngSSdadvRSLdDuNfnf5L3R1qo15BkEmcdfaGB4LToTwWto3XhTEvjuCZlJBdF
K4Wi3qm7/Gn2A9LV3T9wFBKzsHNH+hJSvOENyZTnrVv+tQky/tPCUwBOI1+bGgRI
luGXpnlXezc3iJwr2rG7qkCP5H3a4oIgOhJHMKnpLcToChmqbCs5hxorKPQ8Q2C5
RW6FwdlI+DD67jJ9Pt95OG38NlefewplSNOKuiwwJV0XbiVofsFQ+UGJkq8bUZR/
+rt67B1UF8jUvZbkptuZpq3c8AkRZr4UiF2+hh+4ZBqw0Ab3+g9ZkoDQpSLwkwUu
qOBqxwAqXlsxL5X2ALN3Qx736xfg3o5Fezjxcg2MPVDWNBvm6yy4vjfI5biZLavv
QhY8C8QG2dy1zEjZAfyNXiau70JsG+H3d68AFAXjSbFLLDq7v+KqIqEbIDNLoPkG
UtHZ51bnSn2pDU+vMxiHk8UF+EmbpSZsk/GYqZATvOGME73GOkqM7f06ZJHsBwMz
E7Jjrhd67/bLYmr+kVKbe87nv7LIvNqxxEfp8xv24ZQ2s4d0JXyINX1JOrneVgta
XvE8JQW4rETWsIATjxGgv9BUALkNT0sD8sXlVQfLV0IOPwJyxgH90Z0cMJ1dhLap
OzXilIGU4fS9JJDdNN7vrwh+5QV3D/PmNUQnewuGlM2SSXAahL1e0POIVbxzlkJs
H41wlRTmRSyusDzTRdcDb5sBdwLkduNEVXutWHUFckszA9PnSyFRH7cmuYKR1Gu/
td0NQrabj/PYdBtUcfRCcmYLjjTCyKKHB0UWetgAUIyy8qpAw4Shate45gpuo5qq
wTKMFVaMqJC3nJ4lw+oH5dvgKDq1/jLMe452Mrd+yBH+uXRCV6fSRRGFe4tZfqxE
O9eXxw1KRQ5IRX/NkOPrYU+dOXrL0qSdav0OJrID0BM38OJxNMfdQUozZe/yQvvf
/kKYLMryMEzMxLY4OfiVUvsBm40uwbFXYZGQxD6NQZv0EryCyyJzzhWz79X20pzb
K7Dj9zHvXtb6HQFqxpvWc/vJkhCjprrzg1o9UC0mapFY9fSdROIWP+YjLWFhm63w
X0WZogUYwbILByhQjbL2ZF/2v7OP8BWa9BXex5Ndz0pC6BYpGK4XrhswOkINUh0x
CVmcMqjyDp1cNX0ZLl4fY+DxBb/qxXzUoZMWbR6FqwXRpZAmHKIRv6jzUqTBE5jn
wdA7IWMbDeGedWubkz9ySBiWZst/Pvh8R1FnrTsyN3wacvA5WfdBccfLEXN0PEOO
u65zyX7XYakbQhEMHqHbEVPoBzgJ3LcEz6bt7cZN+NB5cgcUvi8w+jkniHUeWof/
AtjHLwlaQqnyQnRCppN9zSnab3oW6jbAoW9y7nfafKBK9dSD0KUu4epOoU93UYlA
Rn1VXhfpEJ8LKToRD2I9RAEIPmwW0xmZ2HyBY8ujjrx/UKbPDbE8B/Z6FJKjSN0b
/IOuw3Wpw8M9mO0ESfYuy1QHysLWeQFAZAvD5bjxNEQb2OpCTfMJ1DxzAAVNUQdN
DhjHxLAbXHmwiwVdexdZa+zzlzPw69fLWTBe/J2x6hrWo1jDzf2hFuGBCRg26z1b
WwgaHESW5O+X0MSsSpLf/m5XV99gz1dsj4N7+ZOtIPcswEMneS2Pma27H/pr3Nxz
XnXlq3AAFJHKTizDcJkDwPEJeXOqC24JXXgktSlIDMdBW1/30zRQfgdxYnqYg2Y5
2eiCsXsAu1VntPeaKKqF2sk5eOBTZ1we2+nf/vTP1BsQdjFEvs0GS50Tlip28VxH
K9iqzISpwVPByIMVRDgD7UHRjwUsFkkr8uA0aqhgjaWPNMP/PxGFfXJOCnWpcepS
XRz58DPfcxSs33SmuUjzz3ZN6VOja2KZHzbXBJvccc14MrwSxxum5EiBs/olfVS/
xdVoV6BQX9UIFisD2BeGFUd/cR7ldS8i1hH1ZyLxaJu1bv/hzBYHczm6qI0FrNxR
bPSFIrsytoNltbsElG5AtlPjJhZlZsScTsskUQ2EP0FFSdpJbJfXT+z6Br4elwOY
K5p3fGGPNEGs4Rck1LljNUA+RJerWjxKgJ2qoctQdkRWOJB4CuobLiCD2/aD5I2l
ovkZGPV2YaPVSGe95sbzZ4gIP1DqKbWgv4/J7a9BqL69FPJtaGrIbhXgkcavnB4y
JXS5TYN7hg4Gy6nrh1+MEeI+iPWoFOVkX5efZ6fq1ap9G9xgGBHFXBtSdA/3BN/F
qwHiUBJTvQjaZ6WalD39aef0tO0U7jypPaGH/l8ma4UsxVNtYbthspnVRkCF6FXl
CdCeplX3sRQ9WyNW7XkdSFjtkrw7KxuxjIuZeJ7xI+vKAx/rgZHyMExOtaXZ+mBs
BZyIkAH7c7NDf+vECilj0h1uHNm/kcc2tirDn6k8VlPYX0OtwDZnbO38OlIr1I0h
VGnDMcm7qD6Uuey9rTJoJpVow6fhZEqL8cl7LeKj/2TGrG1U6WALvcCH1/n+GyeP
0AZ9gAV+D0hyDK4tOYt9NfqBdKkp6+kRmMGdFfbE7+OxK6xujoJvMdDSWrWFMC40
nJVBxQPDIMgKOMhIzNMTgadBnLzSjklcd2O3DaXApjFVt6UOFBHmz6iRuA1VDZKM
iQGbP+iAUqxo+nLdmTJE1CTNPlb6wLbhMqHzNnC5fyGAVcE2Q3tPxw+dXXPS0oGF
n44GrX5FkZXOfljmCKvz4ztYjclzxCZVFU62ReQtR8+u/Fv5wwgF8Osj5D202M0X
2cTxA5m97VfHL+pit4VnVUl4jsRdIIm8BjXNP2ynj8N6NxW/isRxJ92/2peiDlTI
PBlWb0E9wLbZcrf5Our1qkdioHLMgCy44aqLfa+4BX1nznX6DxQ+7QFTsRQwcPxK
yfzs1h/mmJrGnUfq5DP5XHWaY/CJkqgnu0NcySz7aLvsMIRkPaOf/oVjF79hYgMK
wnRBZIwsaoKJ5EMbLwueQsL8PaBpknW8AzjOw3IfEbs3lXf9C2rpC3cHeOLu3iuC
HjKkDdelSQ4AmF/SK6le5v4YEfcn7i8naIqMFZiQWg4n7MkErK3lrm0ZEy0Nmzt7
3c89eQPHy/B9TcR8RWXOytg1Cd43Ey7/C7n4RIc6PBmqV6vS83oZen6j6qzSefTV
+6/aNyuh7wlwyeXM03vTgMKCLE2drsecIu7urxKKM876TMEvhSFmdPTRgOd7wwFN
Ie9e+ORUJARkH6lVwW+SAzNqOz8wNaTUIXNbTyEOyHiqW9pbhTbQC94kC1O5pSWD
vljXVFrkyhqa0SUcyv7sJaszZF0jBt4LMDicFNuxj0obdq4/lK5Jss+zcMYMHkNH
+qFShMM67i0NunlYkJBUXMnxcrbIL2p+VMj08cF0DzIHiE/b9aEMIpOtluQwVp8S
SX/05iA9R6Zn94gtkIJ/wefF7UWBG7nL23vyTN146ZaEyCwsW+QPZcEbN2j5u8X4
1dVIywwOe4UWkzEAFRMcpwtp3+EaCpUL6RHnyI2JqaBmHw1VA4YZcsQqPC0lg74R
1ijZWgqaNQCtCKxQw3noiqF4jGPCGjFzQxAdpZNcynt1Fnuv+eIjlUQ/i1KvlHmG
6V5PAkIwuz1H1S43oZxE4iCqcPrftBLym6Wv5uwyQxF0RynKmSJg5aigYnGiYggk
DJpDjQcciS/uzKEYCI2F9jAr7d298LdqOO6ctpPRzEgnzDnVpIN4RV7ODdPmEZ8Q
ep8eYUgiazsVKP8jTxOsaAALjHOwTMzY2SPNQRYlQhlcoHDQUs8oq7+qqUZQ+GAo
TiLWOv+OB8bleD1Y5tfQBh+TP+BTS6az9C4fmBo+X0cCkgG4RhT8a3YJOVDPEADj
Kh+LKht1NcFy+kbiBRgYUa6LFSB2PnixpNC6teHbG3sXvHs26emW55Fij9nh4Qqp
+rL8ldV/rjOsf3FC0FFq6ux4ZTJcnCLEgnfOf8jFNWo9qKxpeY1g1Jmtn7HrBWsD
xb9tYI1v/XjwOq3pjA4K6aNa1FkROjtEQiGk6I1qcTeWRP4GlC9LTXZrWSuTpXfR
MYQ3p83s4O+3z6yBiuk4lCBoKn+FJWGRBKzZpWA8vtsVO2r2bicrDCeXhO/ksvMC
EZH5o6vVa4Ic+7UeniDX5wamzqmDbQL8DSXky2sc4auv0SAWt1hyy3+ZAAF/TB+d
ByGPGQdKRX9Ktdym+FDa1nkFtxJM03KXWhhii+a/P1rLxVtrqU77JGi9cT+Oiesv
EFfhkFJsnVMHFn0PN6xu0cGpQPIrOsptryZnJh3HYnoMrpirZ6+g2jZNzJft6mav
SILye/GYUgGkg4gZItr6/41t/kn1C+SAINrUOwrjpXxABkIYIOoBKfkVzPS1g0Pp
z7wvLbfccPpowRHkzfoFFP41fAIsGELrfyL2Zh+6U3eXKzTTjvgHkIKTa0IwDwrS
F52ROlNw6qAEP7KvDEyWA05rPenPIVP+iSVnUqjaEqyXU/5JbRnFmzDqFKjCsgnt
O0elRUEFAkM5TLQ5BlOyGDfjgZUTBWt19oLxzkSx338Fs6ObCMSpKUTMLaO3ICAx
KzVxtQ0LyroBD5qdw2KLJ3T0k2WseqodTeGvLYV4x0+e1basWDo+hz5+G6o/9inY
Z23Xo4BX3L4an/iB5MoblhaXxFWqghgNH6D05uxjZPRZZFRx5usqeFuUqhIGsKTO
nrnpA/vVAElw2VKZ/8S2qVmzJMIvEEwmkCT0TZI91f5+xAqbFusd894jfFwS85XY
gh3NBB+293DgqdFibIenSTLUuLNV9zsVvxUd6MyMJNiqJP29NV2h9WJRlgHg9RSg
iDk1uiiX0rcclg2oehefRw2PJSu9UhlnWVtOxKYKF7O8IMQBYQjIsX09XUC5JKwX
3t7gY6oLr/3FKXqcpwoz8zpapglQpJFMaEwOrzMPRJl67gc7lmbTurfg0XsDibAU
4suSazF7nnbWoOl18jExtyK3IBv+ZXQIPWk+5k0imp5eZh/QxdorZUmEhVs+SWUL
d0zk7RUL2W0SPIno0boqf6ntVAn0KIXBZCak8GsJDW12w9AUJX9/3WDqb6C5NYQN
wBHx3TTfuRCrLf7sJx3Jj7uRu0X83h6VRiym53TI/2RLhIr0YHQAxNAgRT3TP10v
L+miy0iaspDhb8G7zV53ufPOVNrwbacaRIQ00ZPr9ypEEWeSfR00O+a7ofMUOM62
bUUSnvtURYjetge33EMwMsi886T6eLZg/iq/vdJWd7DuLNwJDTH8FvfFm5cu/eSn
shbBhYcQgbTs8V15nXcZfeeWo7IhZcE/QD9vbsUMHFKdc9uqEl5r8Dxe+1LRFIT3
EQJoniXWVCec8AjJT5y8+DyYMpILy7qpct5zGn0tWpgmsrL2grKsHio4q6G5qkAe
1RmSkTb5ekorkt3Qb0ohLQzWUj+Je2Fq6ZtvxhySjnm+MNYwB1aWNPOYYuIBzu7Y
0b0nHvsCuoZP03aOIOMnuVgpb8J7522X8DU1Z2GCTE9c4C8J+Wu5PES/a7zmhhmb
bfgC4e8xAQuSagsQ5TAMRmjH6Z85ON5l8DyiwuIMzQYNqu0Gc5sa/1OhMfbNh3ef
aCehRN/7Jmcn3GaggYPh/KNaaHOdKOCdr7TzEosNryigkgSenKH66fvVHmjkQHwH
cJwsHy9txjtCi86nuQxaRP/FbswXVHv+fJsxJNpG83U0aIn4KMX5o6JVeNMuf1r2
tgeO9oQhAli9sMPrBdwLFFkbiJwwBEXgkSDtnkFiMJocBQxjmhkwfWKkIka3M1x2
mX+e76WqVVB+Z15am+lW9m5A7juLNjzmhoHv+OHToIhezUXu16DsTtje+quZ21Ku
HRdtVGfNl1BiNvkllr2faaclXWnKXy59q+eDlEymk3/CoUiGyScF8gr3bhWn8P/G
9opeTQSHQvS6nHW5pRljK6w7oUURDmEYJQW8jmlAWZ7Bu0GWeikq90GXUQZsayDO
KrbutjVU3VIlM3dlN/C2sFT4vj7/PdknmNBpG02wa+6dXWEH7CiS/dhCrjSjrR6O
MJMHdZaRQ7G6EcHT/+hX45U+3h9MZ56Qj01Ibw8LzTRU1tOXjHi9d2HsQmNbAB0y
fgmLv8Jb3TW5QNc+dNpNshBlwIVZ84wyqQZWVezz7W27jzAQslXpvu0pAzhNEee9
GguKXhgPtvOMVDgsf/zdzAftAIocQ83B22uLRq52NfoNxJ2J81uskS+z6z0ll79/
nZScQPl75xZveSlxjhrg74kRUrHiCqjxAxhmFMw0AHATsw0N/zmA/kEujqVdgAnC
fsmL0cxQ7NYNa5nmtMj//rCNXnewdwCytTW+aA8EhoyDmShrDzW9fvbrTdx9r4Os
j+/+1elJ66oHyfRboT2Myek/mVsMkYbljie/EDsGBflvvOyhSDMDTAg6KE4oBRX6
ExuL6SZdG6HBG4YXFstDf55P9RHsufugmGxsIroPNLDlxwBBWYyKXfL6vDFS8/a1
V3zUg8X5QcrtSkqQhg0obclBqBWhwH1EASvH9Fn0Eu2lNfJy/gFKrFF188vw/bRP
qhoDi6Vdx4/w679CrVHJZPiPeETugf+9PCn6AyjRgt6c9b6myPDJG4a7SxNjZ68C
l+hODpWYhkfSDqZUIV/j4UL8LZ0NCq8mchbqAhuOsnMTCCv/B9vXxjqNTuMhcPAp
6S8fFDu3ohwuzzB86S8iTxkNUytXkxfvpvFPw6stDbHORgFGAEW5lBXcF/ptDtpD
9dg/U5Llhfg2/jTz0RiblN9I45gqPkZ+veaO1fpywq8/U3EvtGX24NslT1YLot7J
UNnnHdOGd2uEigYecjGke6oKbtQryHK5JZDG6Zz+dPCNU+i5fRmXa+FxPJ7p2hgg
F0tag7Oe5NlN8h2PO0otE26YP0d3RUgKfRVblQ//FaO0a3N+ibh++tcXu9+D7G62
Ecn/Am7bZVUkcM0reVqRfenGWsQyaJMkCeSNkl/TwJvqZra1u7LPxiRWK2Kf1iXf
kJt/uBs2ENWZ1DH6SeBXKPu7ndyQDC14LpP4Jx5W81fa/n1g0ElwAkYbZA+rwspa
h2e5GJfZM1Xra0lXXIVtkhgLLQUdDbvPvUgUY87SmcSsut7UOWNcNyet6i0VTBvK
PDNSsLNDqcS8vkfBxqxlds0WkXkUSEBzHcM7loSY/0tCd/on1znlGgEP2/VX/auD
MzFpq69LSEQiok86eRY6phbF/yyCnS+3/GIIuQSoIWnq61zoAxf6ZnD6VesDeyjm
kaZEuGGHKFnoE6ig7W2gpqoU9q7/499aio2CH0iIk3rDuRlgD4aQ5cXFfs3gvG7d
WlN17m8+cwZdvdh2fmBqcmBVuUF6MaQCekcDr2pf1Dxy9MvUoFD/fnUqO+cPnxZD
7aqb221ygyXyATgv09ElWGkeKv05jcJ20i5d8g8c4cP/lD7oj25Ft+4O/FyzIf8p
ORIzIyuGGZHC0CHaZuQmWSMYpsHLnntyJbFwdG28RkJw+EUnUT71imffXozhmufz
lxD8Ieapefo0t/i2RV7SXEYYaJkltqL/OnO2Vw/O5mV/+mbvoIyDCpk4f45HrbrX
mipO+NIy4i6DrIYnPSP1rdX3Ptvi/xek7deKsf5gtRQydJ0HSW7RRZBg7M9f3gHb
H9vqJ2rna+2YA3SSeA5cyC+huq/9/U5Wq0hS9LrU27TI50XBBuSXGyjSm3L5qm/l
6+8GWn8BuTsFW+IMKJf+Z5lLUnBFvwfohlwPRUUjyGlP9nz5VMqgpF0Gj4pUkLbd
itUqohwl2pWnFwPLwdd3+JQ8i3hxgBPpN+xcxSXYaPE07pH4DG7FCFDzN+DPcFQV
U35g0ud1eGJ6ky7aQ0/jAikwP8qmYnRiJ0y02oKbGhhjnuH55aoni/ty25QXLSPC
YxGUgcH9/QMZ5efRJrdCff+5dsUCj/lgDPpZxgfEFszAjXLeSwkAlaMW8ezUPHlZ
lN5AT4QXtOFdXWMzK8jKGI3vKuhsQLEcXaoYFjrainjrladQjFVJGB/fDOYs5YkA
P/FeLhCxwiV52yNi4aXG0cXVNRSHXYdzYzA0MrhhFTFFRUM6V1nX8OG3XjmZRG6p
Ao7NTWqMCHxf9LXO5yeb7CkX6zq60ocbrXuKBq36FP45Ezd/QzS+Xc0DeqBaj+g7
bn5Rrvv5Oesd4/imHbUIz7bynYeFGIqRe8Bhx2esNrgCnBLdDVdCcUPNdJwtCekS
CrgcjP8MXIKAuuhtTn4C8MVXl7JsIAkcqL8C4o3L/QokMWRJJV/z/6ej0gMsCsmi
vtJVuWWhy69+qtF21bGdesxABNxtTRCWnpxp5jDa6g2jzqLaKp/amYooikB15I/p
JvznElHdQ5AgkYHNp8bj+xYNxVboghljnTi9hA4KUc934727oBJeAiQ75EjAxaiy
ekCokVILbCHX9qhQaZowjyZiXyRSOuyl79/O9eBhBolzC/Ht4fOTy+400am5Asbn
SBD48yRfS2oRnET6WYycxad6ZL6Qr4mBZWJ0PkySyAmWBX6EBpM99lMKM1YA2HJP
k8kOoPq9QmEWPKqlu+gjF/Z6PzcoJldiVKshSR0cNWtRYJJEogkXL5ksuwIBJrT6
QlkW2/yMHcAi9mlaZMFwEHYmD7aMK8zvMhoga/uIX2x0D/yfdkMBhdacdkEFYkSf
cmnkvayq45daRYnkGHkfeD/jfbzI6olC0p/2Kf7gB00lIUr6vITbBBFsOThUWdiB
mbKfSPmQ7oXaAKYaXbdNOLkbEJCKXkjHWVNjDkJICDh1z7N503wY+8vgqXlio5wd
rsioNzM0S8ioFgt+Wa9XFrqdipVt3ucI2BL08t7KFFzWcJHT+h1d9FuAsFh/VOwW
haq82iMmILQpDqMztqv2j3Hib9YaLBH+Hugz+nbQprve6YXBg2kncRALxldJ9ChX
opLU9ebsUJwKBloHz3atpHOiQC0vNeItQx6VrMiUHnUHHIbbL6k26coVG/P/amag
ZkRgRUIaJs090UHbqV/oLAx6IqBGtGFnKb1/xCPKPm29M2zpCl2IsVK2MUldQFoF
hhbQDxEpvuSRLyIKiDKDUjy3vj8nNrkTFj3y4KHTdd2Fm+GlXrBNS03UMqDdxhi0
aAvLtF/nWEJ4J0gtoNtyonUvp7+Lvw7TrRfU+vdiDZ3Zg3HzXBiX31PKwNe1XUCS
7HjRETDLmY45HHe4gffLKNrJxIwgkVv1j4/9GDGGQdl/PfDka8K0JyN8WixvafaT
OTt5KFxMfFIaiEP9A38lzTmlnyi0w+fQlQ+CMUE4K32OUUjYEsKZcgO9VSdXXmIG
yzqCl/LI6AGhS07aMrVdKQq42JMwI071MBtqjakcUHfIhWIakL4baL57MdkX+NzF
2LF/ol/EyiGOlZIDfyvnlD+zsfbB1yKLFrg1VPOx2r8GQtkq5MGfZtIiW8kOpf38
MHuNNKWo3ca2S4bVyhU9ku4st4S3lhvtY2JrS2hDYLruhNHNxBpABY/+pckx6Xni
U2s/ZzCNXIhpdg0aGGkbHwZGieOxwKeava/sjFfRyJ+zlr6hr8r+lsyC9snlR1UU
s/3kNPNWSP85+mr+MutHpkWtVw5PICd9V4sESCmhHlCQ48xsPlnvos50bxWIDokA
YXVmi6Qg7iHzqI7HcTtjsX5KY9eHsFk7onICrt3evuhv5i1yUGBCis3VQ4XF6x8z
0feGWU4kQpBYF1E1Y1bBcndWrmtX+2I0ooH2r3+5RZsKbjhS5TN5A7Wx4VEAsviz
qnb7SeskDrZ4INa6vl+KE5IKshvi5AmPFncmGHRRGgguMSptEg0IV/ZPnfqTIrPq
zX+kDJJU04CsL3Z7sC2NbjQzLzAp/JVMX0jMe7GZyhIKh6mp/RACmdXYtvajs8Bg
Gdv/yXSP/uhzvxDLyshMypXpe8SIA9iIzPQm/5OZcT9eibEdXfn1lzoAJeBul0G9
hB1NvTpOdLf6N97vVjcJWdDdoqGr/GcR9kwgM4fuC4xyds51d84cWIiBc5jl3rFS
90W/9pIcWs8JvoYPCAQuPb2ieThAGW2D3MZUMIHJZzRKenQfUSefPl4OMJgIdbk7
NdoXiWvGvWJ8fxgHwKE58Ap2ZA9XIUdhLE8a5bvZblzlbCqEbwiS9s5u6gqSv63j
KuIUzhyBUeOWyjFchKObGZeow814vCx2SD9B3R0M5FRdC57GHCMahGOnm2SqGIS2
GelbKya6lWT0SI5u5kxSt0Njx8JBJPz2bBwSKKMwvODPPNzdcxJjG3HpzcvNp3/x
ECUSOHOzPDaVifqh2BYDnlijsHqko+PWdf7Jsi8ZfqT80p+9wRqml/M56qpAn6XE
15mbINhV1W/LCE0894YbpGO8zP6KoY1hvCzT1nFDykL0WOyVRk5WeuUlrWMBK1QZ
nXsRup3QBpNFp3EBctQNCh7CYD/n+u+dxTS3/jLmp9Fr4WcDf3aHMKV+wcgiqLd3
vvT7cfv21hCN0GiZoJjapSOb/Dey2QJLCzo28bX4FpoZoAbdV+J8ziS+mVWoLBNe
RcAD7JQua7WItc1CyQh6jrXejwr2vQidB0SLUJqUDHBs5BXHY0SxwHFnmkidTcER
7JziQGgdKRWwKin7WbFSeXV9gZhKBWnS/mRmKU+TOc30yViCAl2ZiyL36yVQXfz7
CvZI7uOdg1XOl+pObRABuVBRmxkUJeoGVjP/Lt+MVSm1uJe84qGHp2gSfzt0Vxt2
GMvR/JI8gh+6XbOXJZWtcgfE+hBjw36yFyG/W17WGeS+yvo0KvMWfdFB0Bp/T+vz
/RsKqBZf63Mt7DlzHCMp/spHALs+S5adhXWvqzv+2EwprmxsIZ+Q/dJPSwgTqMf7
EXL0tXpkxA+04oJQP0FA7oQ3ZSSyzbwyxVQgRFcyCDvTzCfK85PG1sVcZZx7Cxer
TMjrm28/JqApKQ1dR6DPYRF7mLgosaAIeAFS9vvnHlxKOmJO9VrBgRRmjsLef4nB
pfRfZUSYLy0po8ZcLJCT2OaDZTMBwvd9xDCsbdMvof1b9tnO14j1j30Up9+R77NB
ivY25DbVCiLHSt8xkoIVAIPjFrx4oTF7hI7NsH9VSZSokF0cz4V5X+XCc/VwKyAe
jKNKR5z2WrP7VgyV/pc5wPl2CiVvvUwXb2Nj9Y4HIjP8tAu9xG3e+/DTthpQLR7e
L2mItXGGjQxNqQLb9ZI+VFbIonXoJSdPWYs04JFelMUybjJQItFQf6/PjXXgo223
dt3jMsksLqeBVOXdihVZk6qjO0XO1l5sspabL+AlMCd7r0DOhDs6mqwnv0YphCZy
Og74nRt+DH9sWlAxCgqkcfbhGQLSCYs9+CMpvSEguws2qNYjQEIaFB9bnRhaBhAi
fS2u/Hv+eIK5dmEjNrsGllnMQVkkEpfhwNnXB6ulSv5Jux3YPaM6tG++7IxhdIR1
G3oodkLl+MSiXfx1tx5z2iINmnpnvQfSNeCK2hXVR+vdOn3HgjW8PokIY24TPEZK
Z+btLnOoPA/OU5SqvzntcS8xCNIg2ZXHblJZGvn6j8OM8XcURAkEFMs+Ss6VZQZC
DHmEtZdHjFsLFRqx2xxMwwGc9IE0OrXDBz350TQW2RnzYOwTesQ+U6twIvwwGdB1
4lsX4sM55H1J4mdvBlj/KlVDdJN5JWY98Ypf2rpvv461/aPGgAzrL8k4KF8yx/xH
rmMuLNFIVDxH76pEgsigZKAfLykxQHhw1usMveHwWooFAtAJdGnCzMgV0uwi7kKW
iFePkPoJGmj6hggpncKl09R5rctoefZoSJKSJefL+gRy6UC1EkTKiHGmpkK+Y/Sn
JJAXxPANmyujdSnJ8Vx4RpAQmlqP/FWzgyNjgvmFE8cjIsSk3ljr7CgQay3VC7wX
lrI0ZuJi7Rcqo0e6guGD4QReDD8v2K7EicmSVNtyravl4GrQOoH22UCL4M4jm/gG
yMup/OapYmfRYa2+49ok6C+/7mJBmKG4J5jWAB6cMrLB/Rxjl5hN8b4JR1Spgl8/
0ZZexdM6Wg0d5CgbfRp4yujFlz2wt1AvvuqqQ7NNZ+wHp3xoiL3bkmUJ/2TWe44u
+5MZy1SYu2ss4gSo3ZXZ3XUQyEwU3Kn9zqmDDbLL/QQeeJ1UYPXcRwX7aLQ9zDeR
ZGn40ejXvPN1lH3Mdq1tjhRi4HFaP9idjG9JwSagASRyBwxca/zII8N/KTU/KuMj
n1VoSf/r4pLlQJZkUMq3uoL6z3BxMorMo8af1QS4a9/v9RrAMjfepfL0DagThDO1
fciuoU2vBOm0U7sZJLQUAG8R/51ptitd4sY7YDSVYwIirj5IXCiBmm8ohpF8RPOK
MbTwJMzWT1wVLSgNzP7sDDSpKq7ke0vN0GT+6lRkU0ajDYa0bggxSNPSRAYnoz2h
/4IFkQLWRFaOgqF+IBlxlDinchn1nm6vMzdzoEurQlqblqpc7aRc/RrAhK5QANut
Ra8kiBI/WHML29xM1BQBSyYCDOvM13o6kYsrY3uMX2c49l5xtcQj4keS9D7ona/T
l4CucyEKXtBs2lag2kjqpVZPe5OtHRK25nx3DrktSiuWuEXfbebRBA/k2H5jcrHT
QJwBx+JQI5ikrhEDk7G5T5dMYba1ZIZw/t+8i1OdY3bBkHJ/tyZtnTms+pHhP9f7
PJ7TFhzEnufDIhanRmY9xpDkQqIcPAxn81brnvuNsoVEOo+2BNTGGuel4Prfvvzt
+toB+kI/oAXI5SAX6qaqn4rEKMA1HQJgwrXW/BJHUMydQfInjMhjh8vcC6ibel3e
l7W/4Rb+9Ej2AojAOOk5JrOwXUt6GU+OLhF2pPcg/qmEfVzlV3q/rGGw8S9n3+9r
+Hlf5useG4DX5qRNzN2kp5zueLEN13qJDqx28tQqk2XdOhuZ72YXxKZvs14PepSh
AAy66Tdb8WHUhdaBu19ish9bwn9NPUeayf7Z7+Ey+/EEEMH0tzIlLK/M0CHYBKNl
aOJ9lKj1RuoRlEvvLsPNwYjX4qFKwoDuRW525YnQVQGhCjfkn9A9BXlxSNTxB6BF
aCJea/pLaMvC4O0TQJYs4XU+S411XL7UP/Ijq1QRRTkte2OhLSoqdPWmo/A4dmN4
DBSzkbMRf/RAbDnBfet4qqOsKnhm8mEN8Fvxmhg/rz26v9vcq9JfWwOL6ciuKiZD
4oR9ISev6TUzn/2xdgw7muxd1vy5W+LYCCAts4seQXV/6HMyJnhKs7hunmA4M6Jm
7TpDkx7GEM068VveB5fcgYTqFf5fGUQtxev0ThBf2wxRRmz6uShANoXhEN6xYxZq
VpENAgQTTfaBWDIBmH/Ty4xTIVBF2MLAESHP8h3E3DU3ROUIEcpYEoyQAtbTLrpz
MpjdsniMMQQf4dlrsp11Zl46x5cczPZRX0//poddejGDypVj8Gm3ex6FFELckzFf
gQM5l22wKwEFfP6K6GfnPw/MaW0wv9WURf3Xk/2ObBG+P4FwnektscH5iXMgbYgD
jpYK0/e4L6nfox1GJNtQOoc6hQcWKakBCOpXeTA0pvt8PiGClEH29BKuVnAUibS3
4QsbiNeK4I9NI4I6mEOwBgHNVM37FwSUBMDTdLYby7Ahnia8L5BEfntBjUHtS6Yt
hMiifhTIiNzTY5V1r+67FQeLqyNL9Y+zX99S/mmqob8N/GGpwRBEYKN3771qSTTV
00v7ip8R9v/4fZXtbAj4K3maDqHvsHK221jeQr4bh89PHG9Y8Uy0FkmEAst1is5u
c82RXdhF/Y9Dkut8EJuZsvPWT3TKRSU9j3Y7kliyVOjKDS7WA0XSb0WJE3zr1hfS
PKf27ikPSAXoxuHJQCNPGFEWUavLXHDEBRr8oGlmrxP1XvChFwuaR1W/cYuoOezZ
fmn6tJzdBsVYuFcct3/9ZKjm+uY2O7xPl4+QK4GzkrAfo0nSlYiwpQMAJ4McCnws
Hb7E7SeAyH29Poz9106rDvpOC373LY7BP2NQlCKJeoU6wL1/NZobsz2OXlGCv+8J
YWFKZdw7FxBb+ugB5jQvp3esKsIlIX5lYHPxESwZpTn/XPSJqH6PXVZyKx28fwEJ
/+bYhcIbRWmEAn0qcCrzZ5enhkIuDELzAJHiVNDKWQzwsbwsSopjJNzy1zv+OTlF
gr3g8YMNqcP5Gj3LuaVM/U2+N5dtIU8Vq9MmG1+BVFrPCoSih3A9W8gjLSMTMaaB
jhcCHfkoCDUeuAykAU1QhZ7kNwZJibQnPPpsQlMv4V/Lmrm/LSSFxB1IDeyXJTtv
Kvg1ZR3FenEbp98qPoOihZtxtx2kYQzApO597eBCyIBa/cd2uGyRkYrm4bPG1278
Hbsyfs1jRvOOfpGs+G/2cjODhe8ZEe0VVc/SdVTa1BDtWi3R9b/DuarmGJlDzAfn
H3h87PZT7zZk6aRF3QFqZ94nhyRnEPZKqyuO7SKVcRnDGCbeEycYnf+17xIIWdw3
sUMRO+DWdM+BsYM3+Fi94PEkDaif2uUHZBhwEgnCTk5N5GW65kaMzhLQX5noH3gD
LY+GFEAX9YNXFthSgaAt715wQduiZz3Dv2LJpSeD/0ECcB13AEPWlEnSnqxGOuGm
1jHJEamRer26DumOuCy7B+9ClZBpt2UMd/uZ0/z7l/YWSqYi1x7pscsmICPou9JQ
Ewp0nLE9Wfygoziavi0Sj6xsmfikKY7V+NR+YsQpQUhFu1u0v6j7TQbBLDcmAN1V
vQ2S1CsorATliVmci4KipvJvuOgAcuzM03gLPuQ0Sax4o91pFiFQe1N89ou+MT0i
Ep5kdht7RYTokpy6eeeO18sPsXYXDCOaK2NtwG/VqTpuWi2AJhMVs4HgwVzZWWhO
gSw0HDMw4SA/beWQOtT6MphkqSE1mUJrulZtYlkGbeKDT3imHKUukoTb55WrYASA
Ozza0Gker/9t+pp1UfpDIGdUEUSVicWUFAfo/jLkQYWzUGfm2KF+bLrMqh4fekJv
5GRA3KstxKEWgXwRFSwi19d6CsrmCRGPPhdaw8YO1dk7RVBo1EXQYQTW66GHEycU
/fNAWU0t6Vkt0hBr1YdlWRQ91XUWWgKHfYcvTSceS5V5dBOytr1DBfacAcydqyxf
rCYOQJpjjGjbYtv014xHu/HvIm1eQ87BrfScYUucbQSetsGCxRSk4x0gG4G6mlRN
QYP4cw8aUG+7E0Pt1AQnEmE/scdBE04fERg7m9BLHtjA3hSOMtubS24AQVF37+35
kLIegKXInpaCg9PLZ2PHNnqmIMYbCJUwfVzAYKodsBLIltdbfReqjFwca6hCF1R8
lkG2fg1IBomSOy1120Gc5MHu0totXrtOhlBfSl5a4ndVw2vxHchFEz5dDm/8Xndz
ILgX+VOySO05LOakS/d6Ws4JwizIPiAoqats0zupuC9wu2o4ABh+56LQJqsblQRm
D8/iA2OvxhPD4eDF3ibQrrC1IMmJEFN6Kawa7xWr2LmWQfKZ0+mQqYiWFWlLm1p9
iA/okO3v5euE0z/lDQT/JC4sg0I7njvave3cM3d9ikOoWt/uzqNxSlzDHH+o4NLu
LkqS3E8xMYIx+dAsmykDnIcrt7gIQK8yGuuI1LBZ7To7OCq5NY1aWLU9/iWpch+Q
5B6QoPNYQLDjyGmArn2DLELd08txSarx+SH4D4HnF7O3iBN2KsLExXE9sphIXxHw
oLWmVDk30VROOM/At4KOcxcP5MZ5U8bBlO+utBms8082Jg8XRdqF4mXxpEmo2JPp
HKT+4YYLisxpwQ7WnXQL6B3zyB3hqcz92RSryiJJ8G1Heu6A81kJ7kYB0jTBEgHz
S9TPdKGOQvDU3Qm8vqWwH35TumaWE9V1SvEaG300fCmlA8M3Vl9OWDXjKqxLEdRs
+usZ/oPa2DcYBPrTzQb5i7EXgjfOGj44bM4C6b1sDN/RGzi7w04wKEwPIUhdbQmZ
WldbRyh435BESRSDooFLnbAEVeOokBOOabNLBHvJgpbJ47kxp8NOMa/Qp2jwMM7a
0kq2TTd5jNkCT3YWjrQ+aEFUq9HikN2ia0yjoC9Sh7umsi1aI5p6ur2iWy1LnfgQ
cAIf5ICwF5ysadc2nXv/pdToEp8PA07ltX3UhllDfK/hapyVe20QVhWnN1tfuxv7
5GCXAkgMWrmpQ8RLnr1ToV7N3ToU++iMB5l9zcNkgNcIkCb7eBgPAJkuMZU19ayo
nwj1qkfhfHKstqYGywCxAghbYEZae8vBHMgAHRrWGpzMrtFt4XPEfZct2/qe40fv
QmwZk3a+Ro4sZB+yOiQaEZAiynqawKmX6m3SiEPo6rmTqRxf34RoDgJt95pW3DA+
r+fmRJBnVg069PROWT1XCde6J2Rz9uhv9khmy9HBo+tqL/vzYJyWefeev8Y4hWPS
mAvlhboHftx4H/M1ovi8mgxZFh7cTZa/vL+WPSVZFaoWw+VL7TwbT0KSezB6Cu/t
ePeKby/sOo4zCgo72ges9ehEVlAwCmtXB0e+e63z2XyOubDmpjpr5gF+7vDmFY4C
cPNLfke99/YFlW6UYdmvjo9klZp1bz6ys7gb9zA2n7hhR78BOjKyCaDWL82Y5nss
u7Xe6LFC25TOR6b9ehhajUJlcGtxixJyMgxD6XHagGd0/qcmWWxFMP0ppmh7vM9Y
gdtfcoSdE99o/eT3wKjZda9lcgRYcIcCBW9iBaASUSunQe2Qm2UP+zgN2Feg8Hyr
mBY9WPFH56jomnUqqApPedzsOeenc5ad5JktiAsQ8Wxe/hQGqVqpxAdUAviuNGdG
H1Cm6oZwMkd5/l/d8ftqbn1dM2BZXXfCVxTXKjt5qN/L5NNYTHUFHK1FLFemQhbT
C6ed4JJ/FEVShssqxHF+smeFm8RT8Kh1ksmuceVo2ILoZ8JYSEmDSyFEOd3lMciu
GzWTwFVoFKLk/F8c6cfmcrbWaenAMh8lrfR/4qKqsn/+dvni3diY0qau3h777cBO
ijliRu8hisTdtcWMT31FgO286Az8l64AeA35MUaNu4F/SKDcTUm0gtoNtagkCmiH
JjgxYyNqAS9fSOMRoFYBvRHJLZ5LYddobAdIti9qUFDLdQ5MmGqzXl9QQGmRi/9O
zAeqZwNzCoRfkH+WdI1Rz2y0h+3Xbet8+7X/0GSWeQeQTNNKAb0GC42lgnMcqS08
oPewo6hqhQhtWBVXj+VqtzsTcZySKxNtVho+0vwD5eUY+/hC9oW7eqmKNCWOaU2V
pFfUbZ4e1c0sOKNpSYUorSwyySi67Vrp03EvKBd0+aVTV41kEhs6neEi/HUpx207
MdrAV8ooGSMffXqP1Y1Gso+zfP3hVKpJXmOULeQTijJz+W2Ph/JUVDGbgwcY7JIQ
Wl4O8zpMM8g6l478BRvg3I0laBS9fyMZIzcDGTliDsknsuceXw89EzblopOGLSyp
e/OMlz6G/zzESu9+Qh44FerCCmgXdWRwZxohhEGlxIARjKBcHumd2vRk2GnzDC6s
Q+tGuMsbW22XmSPA/uG0Eg1s9PjQIVe6UuYS3BIOEXAZ/mUrQPC7kjiq3YtqU6eS
3kNSsfyfKJmExRu/7C0taqvCw3M8QVbhOfAg5Wn8RUnp/h7zlYF0eaXrp607956R
4wgFsWGRn02zBIVFlnIXqBHqklwQcJT9yQtl6IS0ylrWaKWmtnbbkLC9C5QRlrZf
mLsfTyKWXaKwLOnTFfwULkrosA4VNSX6CE7cgzjNOqNrhHua8RkX9j/EQ9ZkSV5X
pHIpszHGnxr4STcH2sFFMifXY6qby7e8P6tuwQ4Vx5idssqHwuWe3nXQt7upd1Ms
iJyyoOK4jRoQu3NWKU/OcxreMp2Fx2vJtfrWemQXUMKqWIkdPX+ZAQRCMLBkfahm
KhqS5/R0vfURIEWFqzdmBthLhQYwwFmJSRqpsPS9PKoUCdqae6S/ZKiCNXWsF+Lo
4oepA5kcvNkSvCHjX8WJyxkm1b31oHsJBfid5N6IPVozrcem+/hjwf2op4n/stqn
tCP5S2+0H34/Di8VxMDvOCZrguXH49zsrpf6OJIiMUiUqKe0O7zfEqMc6Zuplnop
BNg2bw9zoDNJzsiGRuh7RnOv4Sd3WIPeLAlhUiGh41WhGWCbyA9xYRHELCi9u6wo
p37TOVScOoCMpZAhy84fwgQy9PbOTQ5WClryPq8WCk0WGqsJ3eJIXRUH/rpIgMxy
XKT7j/i6nqJjkSjdxdC347EfYCisHKhPlxxjVDI1RQuUuW17TjkxBHQze5OaSWcg
deh3Knul2BWW2z+qEiwfBeAOy0RbrQg8pCG9Fmugu0y0+RFftfwSsAdFRl56aVpw
pGTgJzC9x9J0fyMVTnd4YF6mjl0wAbeLFQYYyliC+g0xzzLSjr0eMCHy3x7ubGd+
29Ofw1sorsMdxon2cpWFejm2CD2prV05sjmHwafOuACmRHeLBBk3k0bIm6J0zYyZ
BW9wG0h6cN9Afaa6X59J9+WCUAPBqCxydH/hhWjA04hwux0yZvDnS6rscNPqWoIu
5GbTIJJx5R6ebizwWzYTuQgaClfVQnIlmaXf2UW2forC+GKDcdL/FoRd5VgvcW/+
LLSbUNLLGgjZY18O7UdizkxqbDFRb7F3s0u7OSDtUY5C3sbPH2uOVduZT8dDpLPM
GzU5D5veGDQgMdpFIwKeT1MiJLQ4Zme2Gfk0Eaoh8xVZ+/4rq0WLT85hLlMvklgp
768vKHpLUHXFywfkSDn23HjcQbJdZrV9JuzRrl6Ul7APmCKwDcFnlcZIicK1X+bU
n978KrCZ6MY1V0L+5MkTh5vTWkpSOMT6uYb/q/OJ3W6qP45E28rwA2i1EYNmSd/J
1slfdEtRzlkWFKJG1QSeS8sqtZeEGxt2MZKFuv5S0nA1yj8RlATqkr2l2CkcwwO9
eQpuftnvJCTYDzIW/YdAdMi3d9kIa8MxthO9VbPpJ9AtZQi3kbMCCkvUdCOwbPI7
eFbjFOoIwc3v0cIzDMOC28HGtznBZ8hSCgNukLkoDKkgnIlZAxP7eMV6pQoDKLQz
6/P5cqZraB4m0t/3XnqJHbge5h+/HfqLHqGb4wosZt0QWcOJMntNKE44lqn/dFm5
Thqzla2XhRC71Xdu6fjOVBBUmgIWZl2XGMOfdyuVi+/z+uT22L1IXoTHvBDEwkkw
H7/Fc4w/TzGXgj17j0QZshRcVqozsqmkhFT//DhAwD67lD/KWbrNg+d1ZL3mRNJV
BzDB9ObNGL/aCscmnaytw2y19A58xBIwHQWxhkXc7LRrxoGg4Ffe9MC9DVA3Jhtu
ItOW+ORcfVte0962JAQsvnSmvlKTUbiHK4AB4uIf33tu9eaMe7L+z2eGsP8vLRV8
nc7VGvTD+3EOi7chOcecgEgw+XJzO60siU0dPHtwV+jo4w7Nf89LqmVA5RlSDCdk
eMujqaQZR3oek+dmNDLaNnCEHQ3SKD03bE/uSyizhhjjEqGBRWNS78fT2bJGSqtG
HNoDuD68Dv25cRS3yHDtZXhQwGEmszpj2FNZQwsgAOord39mr1V/rq8c2JAgi1N2
34JPA3YGeLxHTxjjIt4X2g+Lh6zNYCYE4tF3IY9k6JN6SLHAGn7qluPbp34yinvW
ozfNPgA63DjsIqhlj0iu8Zgf6HbovHMrq1AcPaAwfyX7GcPLk+OEjJ1NvmkybCQG
brZB1+KEoHcOyXrO7yP41k/bjxVhDQxITPa2sa6fbcUcpJX380CvzI+Vs2ELWrF3
vJ2/nJ6Cg2MY/b2qF+kByp1OAmayytvcjzzGNKku8rq5K3HiCkVQB23o83HPDYoe
a2QPSC8xeId8B1xjaNPc+GkTzeOFDvrVbCH0QREhkUf9MSPZMKHP6eBTxdw+762l
Lq3mQPJR8+70QuZfaI59cuOoZFoVCEXi4/y8AeIIEKvV1P9qYYIzDF5Hb9fuWWyM
uwc0fsjfwjbq+AsIbuQ9e0aB2774djKvJAIOOiuLlND2u8sFP2D4rHMKDAF6dPCy
s18MGZeUEQ9yz9PNI8b1JJQZnQmZTMW+HCzi0m/DiWCsPmaS7E1UlwyxSyDYrS94
7Q7VDF+uuayXCzsgRjN0C6tduN8qU/1riM6ta5WRMDgMjp2Mb6Ds5xlf3n1VFmk/
b5AGxqycnIxC9dmDbCad+02L/EC0V8D++VXTt0f5TN41PUkj/AhwKyO+tYiCXMX9
fnCts1CKBy0VEb1hAf5ay7HVEx2AzTFMbEP4BkmR3PBft3g9m4VFrrtFqkpnWliP
SFq8b5QUE5vyyb1JAEKxMf1tIfA02uDAkZJbXRLVmw1xAZWq+uO/jcLpVsXMjJ6E
YQBviTtiL1xMD49S9Nq3GkkuzHZDtq2PB2TTEBQDRspxQh3Aq9qeBhASsXba0I9h
pyr1kg6l0+WKMfdljAkXdoTLJRKiek+UVzpKk5WNPv+KyjGhmW+gqdpxfXZKWd/2
bcqVPwxG2jAtea72S4wWGcvvboD2TZuNYrSd0TjirnsAtRcMzNwcwFZnomA8zpIz
Wsz4MzQefGwC6ui87QBibJ1oNMd4Xr4okU8J10518oJzN7YRirJMktY0wE8uoR0E
rL01fVjp0X5RTEwYwnQc7oo3J8AxxoI/NmEsE+LT6geFT0JPLrEbWD391Gr4ydg1
yGQJ3LPA9miDfAqaX+J2eGVep+oaf/MZvgW6Gu5kRmZZ3pj2JNdB4iKc8LwVicf8
H1Ridu6gIFW1RBCTU4aO3CO+Ah1Y+oO/6u7sNwhaF8A/e16ief3d6+tqIFOKAgtb
nvEBfnjCwCmswt7XhU3trtuvO0ykewu2rwRnmcvc5hndfRJeJBAVYY6Wz4glLTHl
UPFiQqpC4n+C+5n1L5N4e5zLg33IXlFJG7iqsACAFYe0Glxg77lpQDwVPeDOjXKq
ZEU0rwReiKSvx9Etg6RgDNqdvpSYtVyAykrHnNBPg9Bu+bK0U5DVG+oVFps0o5vk
dhT0IaxgvVoXT1AGk1qAwI0pyKLcyQk90m67+h9HCz50jU3OyQ00tzhcLuRPKm7A
3dIjtz9rtD5BcsZox+UvXb6ZBW5Gq+e+6ZiP7fvgVWh2gMxYku10JRj2GoaLDsAT
dH3tv0wO2jBrk2Ual/i0Z2rcHychoiGeo42u6rTxY9UdiDxwjUnR7115wxhs+r9Q
Yw+oNYOa2W+w5D6nU9E1L2mW7c1NUdMn2JNI52huhnDJBKTE1YGNunU1w+lXnZeO
c0a0FEAuACUJKzVa9ukxOyCOIeoGMT68jth3A/lgDxloK+hHVAeC5rWjCcQS7giz
0R7C1eTmHi8ZtHumFkW8LpgejIg7EyPPFjobc5I8jvT749OiyCIUUr2ClfPpYWHX
OjjejglTWG2YTPvbWuTIxrLM9bnxgEEHlv4gfAEYfzFGmSkdSk2xPxki3lGUNkII
Dd0wLSqL8F/e/n7LKu2pLIZSnVFPYC9HvkHr9At92vj+T4ujc2fvroRYcbZvQYM/
MYCd0P6GUr2YMi0UfJSJAR5Krw6zcfsVflZMM2d6PHO8DMT/RnguQfrEclfn/zPv
GNIg04CRQtwmTXcFXoWbim3S1WKA2Fp29u8qGb0Ipy2Q5CQF0aoCjm4yQLfYLcws
IsN0e1Fhm8FQ+V9VvVgdA56s0Cy5NjHe0ONuPFtcor9MELh6TThb09FPMMj7V54c
gnienjvq7sXkQHiu0vzzubNkuxkuC69BJAOGySsXNWlnO/RDt8kmLUbUi6xAMPVi
I0yrHw//xoVXAGGftjq99mQ87Rg1Dy7XSFXMucAdFlRKrGbpBBC4d2Hbud/b1Wxk
v8+dRGmV24ZAOC/BJLjXHuwTpiJyUnMLcdXjRQMU7/5M0QdmfWHKb932TaYTnhXq
lL3PH6VaBkh+bY9L9b37n+ZnOlClB95uXaW5ZUadZrntLp85YGy/AS78UwKocPAT
ETkRR98mx/JSHBw6FrrM7EJNYY2YwhYKcjKVbKZ2eQoGuwBzcRoC4tQrz72KEkmB
kZAsNAZmrsAA8YnuJZP9+RCVbWan945cL8dOIMkFKV/FXGPhLsRD0UQ9vDkE27AW
nMurl5lGk8fXFhjtEpghsOl+2HUwMLm8BaHgrvoFAQ8NY0dFrW6lc3q8HoZzy5p+
hu3wD0AcIEHW8sYRRM8q+7u4LBq+3b/voUBGZlKlcl2P4KCwzaCyBMSp1smUkcbj
K673MOuoansHhfetoJjOtoljhJt8skYl0scUP6b4Xv4Y7j6U3kYf9OLlCwVJ/mLm
Tl7GZ2DsOGf+DrfnFvLp0Q5Fml5oR7O5PBmO9+tXyTl/558t6bLuDADZpxIFVvrO
MMbN2wXfKJ0H9TYvxmHFEymFr8PgmLWK4jLalec5E8a0RpBRsxVA8ZvVU1tu5PzX
QAjvA102RvbtOVkINz4c9eqYlY92pTxp0JuXbq/1ts5D2vS7LtakOqFIw85vZHyJ
pcVcuPNxC0V/OhCkRVYv2CW2t/skJ+iDGaNpgN2MO7qthtUe1M/Vi5Mt93sOLM+R
mKCRxavB95EVY46hkc7lfOzi3uqC0YeTtbPPcJVSIm5HVKWwGCinjX3AcrVlbv/A
41xqJZxYKMmbStO7ybuUM7SG3s08J5lLQv8fCoqVUPseCvRao2mOr5xJIiiyWuDx
3MmGr1Av7gJ0yTFMc89ZfYXQ7sNlrFmxHZvKZ/godv3pGDDzl0++hw9sYYPiJAGh
yo21tlLPvIvHPeRQ0VtrzmP3aITTlE9GTXAtGz5Gq1KpX+tjE364gU2gRIwwbyQA
TZ5nL6fZrZFT+qc9mE8H8LGYYSiIP2+SJ98KhjKa+vwxBYV8IRJeTiK2gAvReRlY
IpCKx/ZIRm/7qf8Z9OUKjlnXZZKvHJZEaaIfy08gLYTIjx7SnrxESJ05MXTGUDkN
YeKjuGyKweYbvzlaBQ2ekhengoE2RDRq3QuaIDFaEYb21rOSJMLZLDqZ3MFcqBVB
8o0/e7gcMSkHPF1pTpK2QtBEKDZ+Y+smfAdFksdn1kxdYgSuvOLAwv/8g2CHp21N
W1zAFW+l7s7SljUlK34V+MwwRa3uLtAFGkW2M1yg7aIGyY1/3fp+sKUMPRwjSyge
+xmEuFP5idDiWYHePTBbB4TDa7j8+aMWg7+DMSSOrzW2XKh+IepTcmnRRmRRwP/a
VPk0F45AJH8A36e3CFxVttFZdNsXFPz1zjR7uBy6Wg6zWackuZhxnS9iWdIYWOs0
8BL1tv1TEM34huaJ8nloayzg57MhSJYGhr/qNXwX1bi7HL/bQJieoc8h8bQV2wcO
/GuzfEdyGYtzsIJO+0FZ3MMzYcmuRgXTDWrX16mP8IqElDFgy5b+HvHoYEo0VD0o
NmMArGHmdIivJG00BxWye1/Uy3b3vfEmtgJfvTLwR3BGlJaDeof2iUsCpwMYMSV0
RRD9PGCZnBKSp1oLmeOOKfQg9pHk0/phJx6W1pLDU8sxHs7YCn+ucX4Y5/L27kP3
o8QB8/2eC/0zvBbZkU06CyKlUgvdhHjwNEuBB4YSVCWbRhD95uYEQJqBbtW41aPO
oa7Eyr2sxEMK6Z9agPwpkEj8Yd4FKP0VBLnF/LSPw0a4HNDm0oZE6441O1m+lshv
vbl4+dpnmIfulSt2B6/fvPpi0S/2AIQ7YtEJOjR0y3JXBK6KP2Jt5J8gYADufg2B
shQ8Tn096m7jBlp3EiivrD09Niae7OGHIeNbeVjgTA2Tw3vlXm188qAAtrbLnU6T
g3G4M47RA/hC7HoZW3r/nMDjeXbCtBZEw7mN2lo3yNkQG5ERkk0Q04xrWtUEfO2R
lrholmtJk4nICllY8ZprATFCZdPdV1GQA9+XKrXBispB9yrRnQ8pO0jnlTjyhtBS
zL8j0GZw/SGOYC7lG1/40AYtHqbOInw0kSNcHrJCxHLoRoclQx8CE0EoaEJUgCMF
57eC+S+NfpkLhLkNr1WsJNhGA/5qu/Q325OC5B6Ve0sPD6VGPeJQJr0wzw+PAW2K
3G6axTEHRchxP6+PUaWBC5esmRymuRe1TrD54jfzpHevTOPQKv2FlG3Lxpv8Ka87
sjq5QE9sYzJftj/VbCN9CposWQACz4fVoOZXsp71dsGDoKJoMbf/N51a5pR1Fzi3
AysIxksGyY3m+VfFgGDYzA7ZFnsLCXygMnkEoj9PLsJBsYRYRwUNXslz31CJ7OOH
//Kd0U4PnN6962iX7nIa5I9MKpUIXvLcN/27H5+f2FAGW5nDp9N1O3H1CYsmDlSw
vyMaRFDA4b3NNSZ4Sch8F/4mgfQt1daKoRRy/7bts6uqVThSYKRgFhD1CJuadN9j
VJVicbYVJN4RRSCe9TG8P3FYarNEfJO0sh8NdpKCOIr5naVWy7CPe5vHxPBdVQZw
owgeIj7SevM/F/FpH4Vi485c4PdiZyhBGQP6QszSKVDlGvAmNu73QhbFg8Z8nYHs
99eJGnxFUipU5nbk0DRTquIkaeTuV7c0CT38yBVvvkWzdgg1Z9MTc88blsQ2+Z1a
OukQ8Hb591OnS/J1jbJsuikC+b/bJ1WLZLMGSgu3VP2onagwGD1s3e+hiNz9qICX
BKIFPIDo/eueVsuQKl5W90X6sERKa3PZPZsrqYi7rIo/k5+MgXt32BH3UTeTsZXa
Ej25FQNqnjMyOh6h9l8q14DkGUrtHEvd9hKx2Yve1T/0BQSeUrCr9NqEPCtb31D2
5WOGsA8/g96hu5Jj6oZ4LaRvutRXNL7z2nWpwY+2hrosrSQdnKApXiy3aVidl8Nz
nFv8VczA1NIMFYzP6cYOs54nTO7D7ERU90ZtoWm7ywUWW7pEggaEXMW3WimWG51T
fQ7RybshIUgC4ZZxu/8koAjETwlzEmPMhqQVJabxvoIa1tN9BAnSvBBUu7kd6fGL
O69/I2YNEwvui0HwosM8Pr5jH88R5m/scd6grS5vjOKPzb+CWLcIlKTrnQPz1I1a
DN5M7nHgSoUwcRv41s8fib0bcE8DpFtCbfnvwWdhIiMKc34rCV1vGr+JfBL3bO8u
7IDRieLLNw6BbR8O9/2mTDLcwKSScL74EmR8QR9HAm5TUe1xQl+Wx5reef8eLbMS
d/QlpHPtqWjaGLgiytHPy1QBGrdApqIPvacK/YuF7l8NUIwQnwEIqfoBOECp4wz7
+jAIX2S4wllwOZ5xF3k2cf93NdJChJ/j4Prr5skeJIQFu4FcIZE9cdXuRYlD3U+s
yFagy29tZcRZvxj1Na8ZCPnsI7WWwh0YDbkbS+oCjxpfM1uDAeR2lUvjm9aKoDYy
lu348yOuoAeFHh9GiqR55yEzXgAec7pn+sA6Z8D7sCW0I87cm4SNY/QabYTvdNz4
/GZrWVVGLilgSMtSh02f/ectmyDgSJAsJ1Ix1ckVLKH5n4Aihtco4VoJSL5J5xdU
BNTs2MlCY2O1MGC6KoNf+Qj7wpZyP4EuPxQ86eSj+rePRPi+jCTPpxT1Bqe5en0W
NYVADJw7ROpkCgdqvtssscKmiE2ROZoETdHkKDhtJ95c+J7CguKMVi2y4rP0QDSr
ECJSohd0/HEyY5/R3J5GVo8YSBZp0vpM4vKMsf8ASu3fS9n6smNmJTfMbW5iQLT+
tjNaAQPIJYy7FUZndz5ekxubOJBvgVP8bebcR4ji5IYbW+/sDt0dwHyhBQJHCGi5
VYbwbwJzPtEU84igl+evXyXPgqKVZ+S+0VvcO6tScazJIIzYsl2CXkkxEyxU2hVY
J8O2Kk2g2AwqhJg5NdMaevEnIUR7xJy/sJCk1Vj06WsrwCXCjLGky2vCn7RXkG8E
48zmRSgNnmNCtkmzcvYaOp6OkmYqKP/UcTs/4IpaVZP1Y2Du3/M80XttI2RmosFz
7NpFbHb3EEq7QkKp+jymhp6c77GROMsLOuTiQvDuLk/NeGmvtggM/YeasfpGKqgh
7TD2heEBJqJVpYXiTjeTuwZXqIW+nJKgCiH9m3FJPUsq2cwffBT8y5qBwsCdI8yG
mD90vtybz/qesXpw66UobEsXXQNj76dTBlx3nR1b/pooAQSEPwWpTC7DeWtPVLu0
kiKCMBkquucF1sYnp0oCmHEDFLRgCto6l15ReuF4Wt2JRult69RmdvyKQ/z1O3/G
WL1H5Bx2tOz2RMpeGGC1Vz6ghh2/SM+jCBAmJHVNx1BbeflQvuP1IfVIOVJqLxrk
HD0nqc25sbUWmaDuys8QFpIBwn9SQVqHXJhbGaVU6mVV46xz2okp7UbQPuPs7cBy
DMxMZaHrycJK1v1VzVcmWN8Un1Hulw32BM7JAm4/8+mOEj9qFYKQvidLV1654pWB
7gmFkkTSaH4dRpWHuUrdZW8ffhc+2ZM53Y+TzaHKz8UmTFP8bkKljm1cSVF5n7FJ
DXIFw52PN4wDlwyNjhfUrrIV8ITZ5E0NUnPFq1gMcIArx6OaIRig8SCXRH+lfFDn
LsGB4XBmcEIrdtM0M0to0sWKPnuPYAHrIB0/A387GL2RzYCvQkOVrzn87YG0I8FV
wiKH9G+V3iWtj2MdQJA2iKXLU7Octf+ENJGxmK3k21S1oguP1BD8JhCk3AX4g0c5
tYIGSAR6RT88ckRBD4W4DFX+/j8QvbwPden+uYiKhRetzJjzy5nv5ui5/P6fr7mj
tUA7rvYCFY13y735UcCSW9gA5YK+OTJS+CQ2QDrx94yB4e8cH5WMfbhy31uy2abB
qVs9weCpDNFNYyJMc5JE5aTtwC/VlrAxDWLz9QrTmxCNYtZpXHcS2OL0jWaKZFNb
1LyskP6aDEjmLT/hIOIDi/4z9hmKMiQFcXTLHe/4QoGaLeVfzuYNloHgeNQaZCXb
1tp3gmY70O4FmPLVnE+qYLcn85saIN75ctd7Ucvc+sYSXpm8boLr/Ul3Kec/1VGF
JZmAdjJL02F3iJkFrxROYGXBzaU1rqR86887zI8zqDu3Kpj28RGtdzxiZ5EP5Mx1
s7SBZTIk1tnuJn7606NgBAPJVNfRBFLbYKU60DFAKCD9ddvt6QUCLBjKvvTvu6G0
uGZJGipZYr2DK9rlxMF0j/Tr9q95SJoQceeHpQJRb7Xk/irgrEYPmzFkv5N5pupH
EBKw9FmJKxXn61z4B6+qItZAY8zQslaSy+d/4XuaLBDvmbLNjE6i54+edhZw4gmJ
BltDIycklu7j73rZgg2eVNbktKQpV6lXBMyNwTPnmAj8BuKm1G9VcDhXjllMPxyM
3Z08K63fr8io21aFPNW+LQdemQd4MHVTMiUXTZrfVWdzaQ9tF18zszYw11EPV1hN
Z7+ZsXXK2pCnHpNGjeBiqseDRa4Z3/D9W5xq93mCmJG0OyTLwxGscztvQ6pU8pcn
ZdRdpvYeQFE1jEO2GFZ2i88QOknwRfNVpQo9xjrjn/Vu5aGmV+WE5QFGzvmiLPwB
1OOIOn2fBdWb0FYUTJme507bYsgPUZH7QMLz/m+hJfr/1t/y8bH0E3NGyzNpVN4T
O1J4f5rGouqn3ViEm8s3Y5SQuOGVxNmNzjSrs6ohhCrKmZkirqW1GEf+6O6VhPlr
uC6iWS/v0xJafiGVZtyyRKM5sRTiOrtbcU+0dcCVU9A8qHTNlrrf0nqlotyAPxkE
MldfMnkHRwDs5tM1VtPkxdW6sgqQpklq/Gh5S2gcqpcTm6dwin45mU/XFI1bOLTr
dYWCillk66qvStdXsvIz2qQ7ppV3dqNZnfVI62P1E6/NreYV5EyMd2h7VQEm94YK
bo4Vs03TBh1dutylcqdSxzOqHuXwHjYwCdD5zB1UxkEZ3+3YvwF/vX6vHwgo3pMj
HhNK80qu30H3hZ3FFTVL2nspLuPel2RQoCnN9Cjcwd/e2T8wket3/rxvbOnYy7fM
Sz3efnVcjQIiqY396TXD9b7RS02HEnV0h+6YkDMz4PdQ3cnUYLH+JCHOT5bVc5wB
VJtKU5NFUaCSWc2HvsjQER3adevqRlET1XYhZ+hloXkI5fKJxOGBh43/FxqarY29
7Snk8kaUu8kooECtpLTKz29BPN6D1RJxTZ0QkNRYOAoAM4EYQAOMMzzP4bEf9mio
hV2zWqCFoYw33hejieUHcKNIbV1WEF0+STXyn6fWxse6LvXCCZhW6m+W6OvjNx5B
Ir8f2DwbafUd3KWpCbDw4FGaX+MZ/OosSHKXsAW+U+Awc15fk7jXCyIXXShhWfi8
yAWeu1dnUkbjPAN6vCJxt7HoeYvn7kzIL9K4AK6cDx3aWCKD4OgeEOmyJ5/SOnAc
kDyZVPGJQxZKRAoGODRMrrhIwY2ST3Db0gzQlZuGMikY42jI77TMRtDRNEdplnJO
mw+7iY+Med9Zl7nZ3XSDQU3ZfJ3W2seaJPKM8CMy50FE+C3hjIUWAokeEqEAZzC/
417BuRhvBFiPuMZgHL02xACk/1QPGd8G+deqNi5c9tzvjREUWroNHXnVZezy8/JG
vawVlSOpegcueVU8Lq3zLiXvIePCeD+K42+wTkdxS+qh8j/zj1uFgjtc3r5NPRHz
9SYa+jfjsfz0Hp0nvSomJ7THmru9GxEYc5hO4iJiKYqo6LMpfWcEQPWO4nQE9AZL
dw+FUW7bJaqvwXTPKf8slJa+qz3BSSGaM1WxInT7igixZrv3zkWgn1dHIFq4tNPc
RejAWzoTasyQaIMUGneap6KK985C99p4FgAITaCL5gvxoEsqCxlfVdvIjt8NPuXR
p9qijbVcZ9JlWkUqwGXc6ix6kLq/nAJRGHEUBLV6oZXTvrSEaAby6d6/EFv5FT7w
1FD5p8wvBNGtVPFpLukMjp/a3/KSF89ZZWRGQOPd4PheVAFJjKwWtyLWZW30FT7D
bsVgtmIt2H2d9Moev8Dy16ImikWZvc4wm103J8ugkQngKYa82O8ulLoey4Ub6KQx
20kbUAliJaRZYAbvE0mjHNskttcuO2eSqxZr0QlD7EvddEZHg+vUWbLbEolHDarC
KsOIo2PeWkl54v0OaE2PocpUhrOnPokKgdZQy7/gWI0SEV66D+rspbkgIfS530sL
zr/rjd1+zxmCpoaw+vRjrPnnLk+FtlWnaqL26vUwkGlwDS6ozYEdaQXKwfP+oHEJ
W7Dv/KFv5gEOd+dGRISvn39nRc1ezJ1ZcJEhVDgrNXM7xNphSGgYnYHffLTr6sL5
cCROcN+E5ks0yjZGxShe1u0L1v5IjHdH4O5NI95HZ5i49vuluZQbi6JJy7ftHin3
IhGkuSDU7V+2H/uuCcWWtVNQDmnexaXXZlORFOyuGSgQ+lFCaQsQMnq/mItlMCWi
6LLn2nS668jYMhfcZvaslfOgY7jW4Asc9vSeqcm1jGGOjr+jc3LhBPaHEEiLh3G7
GlfnX/R5jAS5F6WVupEbFD1xPb3HfPF+3I2CX+0K4hLh9AM4ssVs9KF+i7MHVlnX
KoDzgfAOu8QhHIikD/h3Dh2jpWKHwo5sosCDMxn8MUfrLhTfZlXcWpQNpndKxWmR
qHy1ECQwlLfZlQqllUXQ91j8giQlTHvH48PDjFCY1pxiaixISTrVCzmcyi4jNQ6V
kefVTLDUlLHnT5NfHJUVGIOFD8N3nEr5QOfM5RkmA56mJ71u59VxWMt60JZhmMl+
67oGmzGoYzMAJc2fHqR4adffQZE33qQ4ohTD5uiaDbO28GpOf8xN60P9DucCM+Wf
Re2mL028vk/5q/18hZ+6G5XHZHWZ0bjgPmxuS1xDv+E3sr+Oy3bkfJ6WEzQIn+B2
h8qfrTUUZrjpi6aKSFmaev83vNxplwdwAJyYQpbxKmGA6CJnV3P5e60ymgttxn26
FNjXAPZPWMFut+p+I4Srk9F8v5N7Kuku1WVIZfjyAoyTt9CDsxNwdMq7e2SmqjTT
CuIN3eGZOI62qOGRS7n67ZrcPTtiYC4YU1D86uwkoM1zqk6rRAzslUJoRXTYz7Mu
a+gv8rb2cIF4bRYVC4STQiGvbNKg1AUz9Eo9JT6TVurZ6R5l1ks8ZAvmmyG/EAZ2
HbCel0q0N05KciGmKHoTQc9VSKtIafxSKwMaWReMcxoDNfZJi7FdRZpmDmP+4VHl
YQqY/fXxu164MxEGq1W0T0+gc7hd06SX7xaHApJM9BgF3+w1l81qBcZQqLStoFOh
Tb7kjWWQKoFiNFKbMHB8riouw4styIFIOl56hWkvTFIq0cCvGqgOppp3HFhjn01V
wo4TmBt3r5CLEvz0qfJryZa5mr2zm/gPge8RCpzOGNIthrFfCWTWGcOhoF3u6hVX
BawR5XQEGfm+8wJBOxWh/UVdyP8AjuaLEZyIqekS2J/wfDzvr2i/CS5XQzxYc8U8
tKGGt/YxjWdQchjxIDZnkm+/4iANenqjTspbPq5T80oZp+EYlNnyZUFHtB9EY2RQ
n2/P0eaFA/kSjEUoMFpKR34v8n10tNaUUyFUotbmq/TqsZCCemyMmemMMo8Y0Xx5
h+tKhqaNV2XyIKvNk/yYK1nCrpbR7Xe9W7pUDGNzrOWva+Nez+HQs3pWeSvQrVZU
w4smpgmT6ThXbvvAbWwIgfKYrRr6/4ThkrYtge0f5LYr/qCwWROm1EFxpa0oCkeG
QSXl2qlDjN3nm/UA8ovMTyU/FzN0F3v15b1Hb0ieky7BnOKU0dvUOYq/vr8QI41p
/vRYs5YnCVsHHFEJDjr9NmECT1dVsg3kvjgvE7Xh/H5aI6Ia6Fe4j2lKf7UAOLo4
mABi4JOV3Qxu0v7qVouqLc9R/X2xssx4eP0cw9SjBYKltEiwZ6IhTAN+0FKX3Qwn
8Cn1jBHXkAcp4xvHXDd7x3y5VRR9VJKh/UNI2yjdORUdRqYKERIBf6gXsk57pIEK
lkMIt+VbYn7JxNkQNfkj5F0lbwawpoUKOd4tKM7kIl/Jle9L3j8Wv/J4/n9QwB6C
GboI2zaOA+VdgFifQqaNbOjhYK3bDTAD6AenzdGR4glPyV/oQSu669SYJtlcEdLB
jNTneMgy7E33IX4HuaXs/ar5Wn0QKK2oX+uObOsCi1a8Ri1st6C0Tly7zr3emLyG
GmxXui5sNqTWKPmqHyG6S59ZqokIx2ZBoPW1Kb4d+VJlTXhkagXZxQ8u01llWSrr
wxsSPNwRncwdtgY7/VSHDdEMCD74WGDmGMg/3qQdF3J2mwz9ATePEgT8RlxEW8Kk
n+NJ9i3xqG/TvDyAusnTfEs2uhT3BNWjcRG3DnjBQcP+o8lrJUGHCUiHwBfaszgR
TwEzkXJwSRBQjkadj1FKZqA4UxFdnxC7LeJqt/HvFSu6WWdMMBixngnsqKhlO+Q6
WJKmDEWi1QcreOchYi74+8lIeE2/4WXX7kRBR9DX9jyenAxjxWdszCoEBe3nHwRH
y0tdtRIIj9RSG3rVpWQ4xw3BI+EFMEo8gxNz8yjEM/1/wUFgsv/71SWffs8s8kAm
MBuBGz/2lW7iVJ/LI0AjKS8nDasq1zTgAOCQEtTE5/KyS1IL2LGbiRaVvz8aNgT4
sARcOV9ZaXAd8f9I9q+IvByxiQPCoQHjTrAP24jaDIDPRL5lqzil8ckQE2Wo0Tn5
mDhFfDnbF52YnsJBLCoqQkRgIkJmEYtLqG2wA5hk+4jjhuGjTlCv9LJCOTazg9i8
tFX4d+SFPj0dJK8GF1Dm+uUP5sSMsOItbMqNg+E6bgt5dBuRm+5V8yD3ly0jwA9K
XIwJQfn70yfLhsbxtayqAqr4E2qnTc0jl8A8TT/POjdKMk1ePoWH/3QQnq/0F0ss
fP3CD71W/I8ejZmBZdXH4nE7AIAvaZn340a8RLjbKUQCuai6PRmZBpaikRFPhuoB
Vi0YPsfQCjeT2CuIiIxuhKixHOML59eTBMdpJJNrukR0kNdX3LG8tnNULj21uheU
VwmSXu3hxd4R8P8HwcF29B28IDC7O79Jx0A7N5aSSsw4PaHkGmOEdwOWZHQDqBN6
PO1Pn02hCjK4nHIMmx4EtXCF9hHn0tfE/+HozBg9hD8EVqmEDK5a9/Ge6Jyi0Zfr
FtL47ajIjqHmOVyn6mEeJeMsBRmDUaFc8H5mCUCV9J9wIXU3p4kNR6sVEjVhAqP1
knm03W5iJDIv7zuIeoh50syR8Ke3YsW58tcJDoUCF9zCErR2uwS8UM+QTiIvmL43
Y28xDyXdnsxwwboVyr6jeOwJqFaO4NTsnNDQ+UDVWJZRh0w3wnTKWLM4p65K78U5
EAa0whjsUOHoCCdO9b1BcVmLQhgNaKaMhABiqU8K/wf0QT0boClSAqNW9jJNlEfk
GgUvjxYwYg+2Zvjs9V3GOipLWU11Ijk2GeIIlmMzSjWtxLVZIiJFLuyr47ixYPsP
+znXnNDFtAqj6kxH3V4TdQvvpoZ53iti6XAaivuvjpWX+c2ZDaNgTJIc50LN65Xv
4xz4G4Nhj2DL0cxRa+qdaNCpXHW9nkYo8APgvDIWxM79iahshIIoGwN6WGfrGP4K
3aas2KL4duTvBSJ7WQo1NsT2bbMhnMyplTBpbKgYy+bk2h7jUqEXs8mB4jZVIwWT
Q2gCxkvHcvBIhIMhgrDTbZLAQ4TrN3pcaOZIfavpvkEG8gNLTTI9OMIjmu7mlEKp
BRoD11wXmvbUolm/AE69vWUGPbW+7u5OwlpUb2hFhgT1yL+dS81aPYlFcAsbMIed
CTjFwBdaWsIwd5XzOYamP6DR6GnnUWdSwK5t439YWQvEh+YcUkWsCsz72Ye9Cdq/
iGylwiqvDxuOEpYdAvMu8U1sHZus8wlAm6+V+qab66i/t6S0qaiqVUggyY0kMQT7
N0Tzt6AIg2P6T2z61Rxih0O7gUlpJKQ047/HgNJWAiRtDlXIJ2/ej+s1QpOYEH6w
VDHao45iACa4ZEV159Jbc4A8wOH9lVs0WYmyH34aPTKzZZ8L3iCqJChTeFN71d7+
0oAp60HuBf04naF/uDUgQhHBMEm6Orco+nPM0u05nJBcvfau2/hT9S1CyUVGh9cj
NiC09sjLycvi2spMnCgJD6Zu8pAcAOVCiMR5q+MJTUJZScvX4H09/bmxBwHWflAI
OTZOUdkk0Rt+GfpUSQzfOSXiFDMfl1BUyTBRStxf3jfCQdQbvxH8SKUA7dOeZWFM
zOCt7FKAVz3KaLDmNYJA83X7vFvMXn6Is+eKS5umN79z/QxjwGuBRGHnwWRA3y2B
7Touq+JnumRplaaL1Ur4GR+2y+jRjdteLRxreUwmOFfP1uTwu943Hhc0sWpjxlTO
VYYH6hNZQOhityL58ieJNMaD2rKWSQFLLfQOEOe7xugruE/2kr4cFlJcvrTjE88j
E0wAmWbByoYD+v5pI9I0Z7Mb5Yqjo/8abTk9w9DjiRtn+EL+aZ6XLhL0k7vRCPSl
B0Z/N31/izPmBh58adZclxVikX51G/r+pbt+NSAgoAz9w6VKP6zoxiuliqcgipOv
B40c3ju4sOWKa4XNzn6OXvyq/KTI1OxDHKAV9sEEuPftDkwJG/Wuc77+Zz6xofyE
FfItbcbcB+U3xgiGPazMq3wdyaqxfMCJGI3ffvfC+i5Rs4pK0zNMVP9bdRl4d4Ny
p5+580c/8wYTKMC5Ket76v9xlKeHLEQBIDLpnuzhSDwWmv6K7SyXBryaG29h3SbE
xTGJidxFJcAgcNt+HkGIWB3Ty5dyvUObl1LzqctiV+0sYOxSMqS956dvbvdNWyfY
NurNs2LfjhMFO/0QA7JGFfRpJ/ofm10VZBYYfIToo3BArUE3wiM6uJr1qxrbpfRy
w6EJrxxIVKmJSedF5CoHZpNcTMCbDIoZD5pyRR5atkR5FV5dd78/bQhc2ItT8kkF
W8PQdE/gibSrRQDV9lJeG6F12P3n0wAvdGsPXfwTORSlR7MR71DW2rrIFbpLAPTc
4roWuawzkZ5ZPPwx2u8F6QuYhUlWV29mdzS3FsU1ORmLTPIMAQSkf6yAI3nol/Rl
uSupSjC7AzPdQXMX1jG8Oj7WaPEvmquld6M1lvGQkkvxpSxPL+YeuLTwR2syqGeO
4szIAMxiMZZr2PKBTyLwZp8lXIBV1Zw9ZZQZjSxTZ5dn9E4O76TsM1isxLPfcZyZ
yfGMdemgEf17aV8k8kHC8b4CSXwiSYZL5l2vadFFmdcnRKquYMW22rBeojb/3yBO
q5Md+STAQYu8JF8rLmKHjDin393v5geHTRkmNBIz2uhQNN4FB2LVmwMEMibh77uT
h4k0RGSv/I3UgZT7ITGlwtqlBV4tYO6DjJ3Xc96oVdi3zYv6ip9g3Pqrn8A1vc5F
0evVdtDnOu33kX66/AZg/GB0MQIqr3/SkvQbS8i6BFhM4evc1lUCt8cxYqCMrXL1
hO7Fsf4qIsvu6BLScQPjJ0jX1RkQcrrAdGHxuKS5Zmmn+q09T2mgEC1fSgTqhFOO
t6UGONW5mMIrOvLwTVSURRrT+fI9YjoZUl+EuuTNZdmaul3+p5bHqkm/jWSh6xPu
+O4bB+YqAPsXT89E7AlsumdK87uHbaSdvjdS2vGQudNjc2xPdB62rHTBsnb+jXfl
b692rnEkMoTuKJFSHmp+pkaBQVdzE7Rtqk3Zb1jW4VECEWi75Hjjm/XGWplYL/eR
/RIHw3MX/VmEieuHC2doJSik+UUwSggfl1pMVfM+Mk7FOWOxqkNadXfGQv2Dlekm
AqT0LZdUvW207ycw5SXCLL5kPPg0g+/RSuhB5c+sLzI0JDMhuZpeRnxamTD+10Qn
PeXXxBfZPHUQ3wSpvvRPNoaSV5Fh4wipuGGzdGCiaCkEYdZKSsS8v4Ib4hvORea9
kNWSZ7L3NORYq44D4AqyPHqGSprlpj4eu+6UXKxsAFrnWc1CE6WyKXVgVF9/QMxd
0uzaTZlz6KW2BPJkgMfkBDiPNXYQHlqWUTvRjPKDbN4X/S4MlpKZETBpUKJKymV6
P8ufAdwM61jRo8ersM0eQtX2Us7597W4RpNsaq1o9/bkU1l9S5gqRBdwl7eKcm7l
ZjGV6Jp8IQa8iC+9ikaLTb77dtoG2mdI1U/iZhaRQGWNcLh/hWlZ7nzHNxToq1ab
nLoS1nisYrSyjRJfvxkhPWJsvRQKP+lkyRPBoUO3fH77Crxr2X0419G5mI2D3LC2
t8G+jEn8bYiM03jriixnTFX5BuOcxbmYQbD4lklNmLWTW5cL56LMhfm7eIQDFc8V
vM6c1aJ6C/pXhIbHt1zf5vvDVGYqsqM7x1HYmFrqI2FdNq4o8JHbf2v76MU8ixfU
U/44BC8cusHlBz9Eyve/6Jr0Ke7IEOXyhw1+rE4to1lHQixxCJYDri1NNqIm4Nqb
2FWss9N2gevyV5zL2iw7u9cLw2texZuwdj238trGAYVSpECzTBMj1WRqus8i65t1
ESmUanGKlUfaZSiOSbPRB8BX7IlYcQfmFnlcO671L1GKfAzofhjYf4EFUI2Re6Pg
ME6aa1h52OItzSUY0a+m3gJ7kxPlhOeEiN+GRa5s+MEJESA7B+8ZvWB2KJVrGy77
ccyp6725piTYka9E8yzgeHO9FMatJedRxR2xiV8WgAPJNXzyO/8C28IgkbJPh6Xk
YZ7fbT6sk6DxIc5BnxpNJ3QTeqA+U7ugfLn9p2pc/kKstX+N53+RqHh8Fjv8NCEi
i/jNA9vhMnLL207pANdK/b+Ta9R6V62Zms+tRhqGeGaKX4tyZbRMCr8RyLW4k+MI
n76ZPyEDw1lPSy2RJVuS63AggiGndfHAjwM/7mI2bvSqgrSveYSOREIl2AjiyRqV
rnSLgk9ItSjB3TZ66yTiQ3Ge8A6ec5Z8Xs0rnPLxcEJd1GdkP4q/4ArtY/jsmOYB
VIHNkhBW0or3LPdNlJRSmtLAm9U5784scHzWyC1jI3+TN7Nt2KXB75CFqBA7yV3W
JoAso6qYHEvprNVuqDcB8zdT45on2fODbitZIGdgPCanBgQg0ok9aihn0txdhtr/
wQyX2SP4UVCX2nCUquR4TfEUAIpjQT8BVn1ZPzLVGc2ChOxGkAyGWHVY1Ycs5cgW
QUVL1iP6EhjZfy/wqUF81JjjIf9dGaH5GgHxX3Y8ZlGsRGDtmSbqJNv8hGciOsJh
7eHGDhTuIkKRbPVJ6oo3WfBLXjraMI0gs4cM9tQypBH9DUk4+KbR27ueRLK1+w0W
rsCQg9+5qqNR/gHOkppQskuRJyyCwtPp5FY3dwA/qUfHp9N12atDUG1EzciDZMRt
jEmW8s67+cjJNPCPCRGyHCZacFv9BQxHcAEd/OILaOSyF+Ugeil/Nt61g/DOSahZ
Q5l7e/2VSDoUZRITK6AzJ8lzefckd2B3kJf9nnCZZ6iyydGGIMfWhAel8vvmHrHv
woMDHEKa9mvfeOwQOyQL2kx8DQ5zjAYCcM9BLkl9wskR4YGOBzC9O53aO1gxkjGw
NqdJjhpXrett6+yhitsmuumdCvMWHmiBuWCgopYhfXj3O/TMzYDmJIIBCDzo1A23
4QxL45ralhtjlrp/uue6+rFurbuBo9fmocdvTkvgx8Zo7QTNkwGOJugw2DTBhTUj
5QSCBhRnYlNoFF3pwgcwxJdn6jVlkB700ej5V6kiQbtKcndGpKFqcqc7s76Qh6ea
yGpgA9vhcwX+K2KwUb6iRSx1k/9IhJm1zP9iifzU4W9jlQyJFohMAqUlDg1tWGap
ENPRasUXPIeFwHIhSu/hHeHNE4ZHFQQh7V/SfKFn7ZIoTc+WK4xvQgg+zq/4G1tF
OX6JBZLWOLF8Ivj0lDcDU/RrN817WUejO8vceI47aANZwJ3ElIuQev1c8roYLw6A
zIo2xxOU4K8vhtM8S6KFZW/UxKF13/w17Sq2K9dLMF6JoqJ2KrtsjySfPmCu8qgD
XlE3QwsHxalQwpONm9jm0j3xZtoNnLYp2elBcwEyEgFTy1863utpSfUR5nB+hcdP
dRUtUUBIOAz5WvFy0DYXK52mh1qbPBG58qFo8ZCj5OAX39nns6U7arRLkZUTFOXx
u3WEIVwAfx3KdcsdqPZrIBN/kSS5PJYo31zzEM2luWwXpzTkcV6L4Y0VqFT9sFf2
OEtT/03gCStDG6bV/vTp0Pj5SRINbHHp+Lbup4u2xNlx3+OXbKi2z7vR3PTDSd9T
sJX+CGkEdsUKW13WOhZ/473k1wX5OpO/HeEaZ+Xa8M9WCP7KstTw3fA7t9MHpRAI
5269q+SIHCUd+fiSIQhHRr/lduVuKowzN4KjKXggjusD5uduwEqeA7vlxGwUlvBX
Xv34BsTUYa5Wj5sKdJ/RCx8Wy2hhxdVnqSIe3fAOs1CTtw2ZJUsytxqD7XVZWHvS
ULKM5Sp9X1IgjBsPoHVzchL1yls9fpw1p8Cn2nBWSxwTfZKAtKFXz2FLYkcJJQn5
tCWwzipVWx8wbG+4vLupV0vD4b21/82Dk8NAsp462fr6+qd56K3rdJMBh3ior5K3
Yyammhzr3Z/xCO0sxn1hOgCjhlrGapU5uH6NC0WlCxCEJnR4yiXDHKhQRCzMos1h
tLgiaSI9zIk9VC1JNkmidzCa5LaUwOTbXCKY56vhvKcjFT4eWJ61v1fS5XH8saY2
ermseRi6gIRYPl00OQE0aE/XQhfyMVdfIRWkM/agdkFDduSnQ9TQTn2ip4Hun5El
+e9VrqgOXy1Zo9+xbUXn/6tK9RHY3TQTShghR/jKsvjAsqDkgE0UsV6ey2RdoS9H
1xCDoKjS8fz70JkvjFLwdxkKLMPcfRw5r6812H3HlxjqUkXuTTAbgbAF+SCpg08t
CwFdQFDK7scb/5+RSBGFJwhIh5EJh3bihzJ7XByUGvqMhyz4QtuZcQ/mUiZP9LoZ
M/istLD/YVMlfys/QEawkQb/4+EpsUFJ1K2MhAV2nq9yUbqgvK6DPR8fmBy6ALHg
LNR7ZynyL7MMF6CRvGptUipaclCIvjgW3FmD73yJQu+fvOFLBTwJ0/apHOkuKAap
TvRbQFMt+mzd8IWOTmgn277/wmscmaos6H6C7GMyp+BG0fxQyWkkZuhnq54mCfmT
WFK+UlUDBS8f8t7GfxG/D7HP/uqyE3ETUgl3XQHLXZvC7Z+Dat5UAuOoBfhw8R/n
Wn9Wi8mK+XNz2j1xi4lR6l8exhGRIgRdtPPvxGqFw68awuRuczKVeMRuoB08v2Zd
lU8WieMDfD6nbF9Is6iESaGmPiq7ULI5xLEL0MDh7o5KvZmDQzii7z1GLo3gkntH
fBOa7BPZZ6UQIOQSM5u3Smw+Kc50V4YCz+oGqvw19Tv7Ak7k7GdDchONQFNyQ9QC
lC0l79bWwDInlNqi2a+bXddMeay0pTLREVV7TJ1oNjXjxvuxvgfFgto6tphVMdRD
Z8lNpFLQQLHMeh44lSAUYyMd10pZJwC89Yh7HpMhyfXDubMuTBgXXulCPnO1C4Hf
zOFQ5b5u8/t9uoTJl1GKua7G+LKXYbd5K5ngYxP7VcF5yDbiuMFN/kD9QTT9t0oz
+u1RQttzLifxV3X3CP9jZtBBLtxzNXtH9ckWCH8SOPv+6/OLfK55emgVYXNev5IR
He3sNRqHC+85LkIDZf7Byvz0GbKiPOy3AGGQZyVfI8rSyB4e9QSqw6UB71uuqKAt
xa9uqNzFTZH16yGSBHp4KPaB05vxRXktHQ+7XYdnTJPDb9OLmKW39LFf4NF7qw6b
zMnYAaZmHGjWu/yPUedet0ObbHA49vVLkRxqokBNBMzngEqdzZStmNLSpeVBIbjh
RCBxH3lGFW1MY9MX4gUnSSXlD7He4BTpJUqgI4tEwHDItAqADQUumdLUW8NTapT5
/f8rdrAeL4OeM5kjWy4TH3NQJcreCL4XyYVAsxiS4B3YQ8+C57LoQfavgjbjoFo1
afK/RoaqAKkV6YNUQJLVVk6BvjOhDExiNNFY0AVO3NA+E6gPLJIyhG5Ox/SUtd8p
aco3Ek4eGyLHZoVgVuTVtLgzskUTXxyaS4B+vt2SL4t5NOCpMj9C2tpuh4e00mQw
kyUUHDcWx/C6oztqXrq1/3T7yx50YwuscBtoaCjO64IaDW4e9dVBDl5GxEYDCwDh
brPDcO42PI6v8HU4gZWeoLzVKtnbVmb+6zxs6lQmpiHQmZ50Ek3NrEeCjLYZUmfr
eZjnY8BtxXghs8Lml5/H13SpwS86sOf+fVVDgWQA178NDa6c/00hokKpoVJ7NCGW
xJ0t/b0W/JXl21nWE0kXGUfMO1s2t5Fv/Cgt6kZ/uO/viPKiUwLUC/qI3CRe9gif
Qxfg9YrPAKqcHk0KoYUgKYpGkle8iEFzmzDQ2Jy5xXD/grznJe+i6h19vD2olPuW
ml8baT57BBxd6juXp8c7+nDGb1w5b9du0rIemryxghRTDioS1fZRNDAU0fRGOreh
uTDbJpyJQ8cuVla81n+NQ2bj9PkqWEfS31q3CpeK/VzbxjMMYL0zHRrsDS5f/djO
eeJP8N8T+NXFXidWVq0VXI3hck3Okc7PnOn6mu9Kxc/7rmygVWFuLy6lV2RSflyu
ADuV6/EY+8YmOloIq3CTFF4VUfTGXVWMIPirDBlQjuE3ESVMmWyUixXasjAU0ENH
IK0HWXCcFNuoD1vnNdUn7MjtcJkMQGsjxF5GyRJb/xGSIoVA2FC991V9HcV6cRcw
baDAP1rTflbwbDUhvnyLnjudb2YuJCr+2mSxiBkh5o+HmtXiCVAHo+MUOUKZ4wL+
bQ04Itoj0KbF9y0J81h/1o6rzQnCpu7lKG4EY82DfGtY4MoRhZiSY03qx5KfEtDK
rREiRfE2Kg+n68nfx/CZQoQdnxYJVXhB6qALI2xc2p2Ch6csKzzOvNsTUNsBUiH8
58gYOqNuv7Fu+J2w/TrM+tmwa0L1hvvXwIVaw+7BI7TR7m335QI5JGHzEz+Q82Fy
oEfu8VTkidbJNwufBS5s4vNEe2fj05E7nmvN5jvolY+nJI1yz/ktwZpDqfWNDAUt
DiAs5KPi6QWIUWHKahccA+AMBomQJ5R7LtmkhwjIJ6GsW00uCnlyrZc+qYxa/pDg
WmPe7O1xkEK9X6rP98tmaJHsDktWAqDjB1cL7vPTxEiblv/TQMeGGbI9SurcmfqD
h7rsedcKmPEKcytfHFjTZSPut5lsmTJT4ALFJ00+LUd9QotPPEAsohzP7C294a8e
C+ONYzIiBFruIJ0ALiWdBT6hhCeZBkyYpq/oLG/u9dgRoO+CpohW7uUApTYdDQyV
o5NsjqjYo4/Cfj5z4F0m/ndUvb8yQJqK+8QxMYwZbuTZ5SqDU6iyKNI/B5OgNZB8
TpaMT77DWB4lUgCwD8L7OGws1GytLN/CKo/sdmTx/1NT61AuiJDyrb4Ug+qc/jwC
STNOxOR1nBuuXqNco8y5733FR13jxa/D1Ii0atD/GQe0Q4eyH5tCb73wDlZMzyfQ
rKNqdUIlUlv0unOIqnYyvXp2yt3oz7fX+a0f+lSKd7DF5TuaMHnybVekAv2bCYtg
73cRkRu8ZKyUKmZBe/UXpkJamYXQIpzSws2nMPe2GYoNoT5EvaGHqdOeTLfaV2fg
1QZU6PXIWapqntl1RMft+3QVy2wVX9Nh4CGkp4IQtWf804flw3Yq5BK3C6xPFJ1d
YkGSVlSG3u2/CG7+48jFnjguC345gSnd6tljZC50ULW49N0KQe1P0Qoh48mo75uC
MCTYk7pE1TIaF5a3wABydEaJA7RcMh7kDlfD12PgS0u32jSDv3IbaBjPo/DvcC7p
XjeMzoO6xINPzjlo34uM7MoFdGHfCbozMV0Ln678WdJCPYeqE5/jLPPh/iLqCjQP
tyu1wr8Vi5KCen5Jk4M4vjhedF7ahyf3vLW5jyinosUhU6jIB+4PdLHyBLZ+wDhD
sdgRrBXugiy/Rioeha7N9ODDP4/kDPPhW2ON4qQAAKwWxvKoinAm/Ke/JnbSENfC
TS8t6NYFaT2jrDADhAJxg2GZwSDruTnh6J6WfbHsQRdqh07zNWoXl6r7SQ1SkF1L
IUnqdZ2SxYI9GbMkKVGgsZAQCE317MY4qqZnd6c5qb9TsLdC6aXNlyLXLSC/9kfs
HG3gI/+1YNgDn/3TdEsnMFvpPg1tUj+SjSbIVk2yf8RWDromaoTzNO2r8dvgeBkj
60ahZNBIUzjZMIStts7zZiPpyUVjS3e6Wy+zu5z59tPih8lFKh1XFQEAcsjSynjB
WP0wvstSV3z5RkVfryNyKGum0u4VxbP3GUpMPJSYiDXkzGb0CXX8bhAUapJhc40k
3vkEj7mRMaD9j7E1BqgX9gxJMcKj9ugFjfD6BKpUJ4OyclnRqjnWiyqS1PoDA4sg
GPOqecOOBc5qLU7p12LhiJe0wTHMe5wtmbh8lk5W4M2Qkd2Pxjdm8Vn4pR3YU1Xb
cUaYQeH/7lWEqoy4Zy1U6rY+VTnOhSz3bv58/lUz0wvVE09VGCxOkk/lIRtMb4DK
xfHw5/NZgDMzZfk916zOORlY6QovlQOQ9j3kLxe0Sj5LD0OwuRK/EuH/303OGJ5V
KJM5CwdFK4ffCNA68/GZs0/QMuJA7IW8vpVUL2DQzOc33WdieqjrbqhgfUT5QfOu
H60TqxkLFKk0xfYuf4gqB/EXpyPGRH0o9uL8t08PYK2WoxTNdQ6BzyYN+KtcswyC
MEC4GUlVqa3zytuHcp2WPO/rXqyGwEhgRb4NGSEroM8VuDYcAuziHOn4fTr8u5wM
5GPl2i8hpU30guLiXMJC/VnP62rsRq2d+h9ZL7xS0IYVhOeSwA4T8XVclNL3v90q
4D1jqnIdgB3TSBX2EmIAyExGw0Pww4sz7GkOF0rkf3b5lviak6sr3GOaL8kS+3Bs
YihIkHyfxD39d0rkg4v3vDGQ7SlOX+SSChDQTyZ1mp6xQYH0/E/W/4/Nh/L5oWQi
jOG3TjGVhHZu556j965XJqaP9Hj3bnKtt9HVYpJA8IH6q9BC6VAyi+ZNo37DAFMu
OdPZ0SpyPYAsF+ZB5B0wweIzoYLrZHS6Y8C/74wEUqB35WseQMV17Z7kAJojKrwj
jvz1bRESGUkjVz/9xLaVkpkMW4m5Ytau2U5UyugjAvqcEo2xR1dHJ1YhQHlalKqg
E6RoP+kT5fzvKr5X6/Njc9oJh0ndjXlH5AncCWSfU/AomRGcW5TFUJb0fboRDAwS
4WutHhC5fwFzP7yPSvNvJjkkSFJ1B8JXXff7Ys1T//b/p2pvl+G+6RieZBBCIGsD
l5T6lF1OfXeAe0kenr1WwoWq9oEhhl4Y5menE3DoF/8yicCUqwO+73fDq3tXThOr
WJK23ZJ8wqMDQcU9TYXPlVr6oNvmFcRWxVglVRttxislv9fZvaEvEycJdaIme5w3
WE/Q1N9i6J1iANkJGfbO+OZXRPj1X5/y8vT+QZcVA/z4FdoYExLWIR5SUcIlFcQr
V37ZmGbskKYyeEcMzJhSPbTOa5qaxjrw/SOrClovxRsYCgQrpVNQaX4HiPYtr10n
iV9sBpZq5zjCDflb/MKYojk7nN3mvYA3WOu3YDHqU/vGnLW520WFzUpbG063TxKJ
KrB8WtMtk4f12PUfCgkSLDN64y5+s/rk5OjlhuSHGtHZLruOfZrn5NrP2wx51CyN
8pSUjB771UmYKwu3DEbYyVQbJx9cZ2BMmUr3KWe1yKVTHOM/L+wZknzuNy8/UzN1
RpCtl1VkVQZd1Bf/SISse6nCQAh0NuHaIvnckjPy4WtTnOiASJ+zMjysy1ePXTVo
baxSzD6YpSmBCPfBiz6FEJXQnM8l2BZRcciwxewBkOCXcY/homYpPi85QMZiXfNo
J1bZzBKQnoFw4llmlgYbwHNdcIOUuJiuyfS6ndW8UEHGK9GFQIauqEGWov2gdqJu
H+tDiPjOo7uvsBAmvBXl71sf+d2bVzZn5NpkaW0r+Xf1OqvWW8EuX+X3NvlGVMS6
qTJzUfZdBd/nwJkeULLiwA7DNN4m9QM2l25lMoN7gNiZoTuQ3ZAj8JUXIDfu1Rft
1UydRsEC/Tq5poDwJGIKp5Sm2wfGUA5nwYojV/5P2+d/g1ST4VEIAVJz2/OV7W/H
JI2UMFIyPhZ1WEmHSco2P+vq5VxBKgs1UGbqSj111lAmN76kd6sXk2y3Y+sIqAhy
b5sRmmnNYhtT0FeHa1m2+J6WW8g48+VAZMiQSZ7HCUXyWBVnurc2DCsPNyXUaLjj
grqAGTauEcOpsAkAmialjdH6yr6vrnaPW8lXdp+avF97JAp2yinEHsI79sndwUvq
m5gQsNLJUDaeuIRzFlpGjdGJGAYcYPL3oxX440tKlpaZHiPzwnZfSH7TJxTZfJvH
PBau+H1somseZjv0BeyI3aoM9OpoNrq0TPvdcg/LY3QVUsd9mwG5GhGKMoDgjpCt
UWS5FeKUbB4FFLRs3D9Wfnf71koVh1zRvgW1WF5mCxCuqj+ttzuPCM6vP4/rbcV2
fzW0kybRdtztq+5JKa7XPKuqRIl+ezutYY2dUZQcti/bRT6UT/VZM8F7gTcJBtnE
SlWiZRvTwOFqu3HrJwH09uIlKyZdOE/QpcK68NDZVMYAM3UcnkvVVoLig/67Xs3U
ALunXU4WnQ5axGeDp0uBijDcukWTQ1YBKMPz8X7zb5dPwpDByeqqC128f8qFbG6d
KjgchcxyFeYWQfvv2BUiwh4pPtb3K+jWIjNR0lJWMm9jszg96Xwz2DgS2CqCChB9
ameUi07qNNryzPezuN68UYhEKnOLfryWNruDdLYY4ROEManTrNlvNfZWp7AEOivw
DgRB4tjFNcpbmLCKPCoPYrZbQbGStNsJVqFNXjtvMU1MKJar1ny5QrZvLwH9+nfP
tH6s5pIfTSGSSNyKAl2dHlJzVp/1MDO2vsDW+oaYmtTVK5ixi4rhepmTAO1mOqTW
8/IvZw00n+Fn5ueACVqVZcz0WYIlfM4EZXVpzSE0K8SiWwDDibPqyVGTLkoHnFNh
WlXmX8S4Wu6XhKHkbovunD8gh3dfEqSm1lraoSsPqdRYGopSRcmlJ0j+97R4FZl5
KoVcRzr/CoMNLUDw6v8xNihwMUSrtTyFLo02dAUH0iIF1q7Ek2dyWOYYqpR5QVWq
Z/1/iXG6bs4H7/WCpplru7kIxlxS5e0INRby3LCQ3NL5UKXYS1pU746ZM2SE3fNE
PWeGWpQ3IjxCLr8PnT6DmlrKNJXKbR77clYbR9pSIlqSUfbN7kM4qqb/ZyRcouaA
+n0ObgIgmWlRc/ZZmwGp4ImsftK8FZL8XP3SL0b6OcJkhkDTk6CcyVEHRl2iLx1l
z5u++bsbruvj2YJq0bVZRYbmEAgX+uYWxO66CjHCxz/8gWhpoCHxRHgmCxhkEAA5
tBQJP1vjW6dkn6YyA8BmwsxCpUOu2r1GVkBrZKvGlGaiTC6RYvFqNIAIhq6k+Pzj
BU7QbnTg3dU3rqKl5wetF4XBH39jdWjhdxyJ1lzPnsjkgwJAwb7PONlsS9mI8pgU
YC7IT2kJoQw6C118f+OJjyswAOgF/eZeFfUcjAwve++/6aQ2fes5OB/+VcUVYUG1
Pgg6J9EUnElbXIWIioPuqKI7S/+rSojor2i6oZY8mS3fGbwaRKfBb5PYw9JX7qyT
HLlMPxXeiBYjDVuMTNm91Vh8JwIMzNIWNk0XttX1QOTwtYCXYcL32XkNT91/GFKp
YIEBAl3T8aryw6b4QXc0g6T2kpM777oEIV9JbaiMwuhXBELoVJtlc4br5ZQjNUsx
Lrk3IcKuytDlF4m9eZ5LN1sUWJJZIkpeMb8YU59OAPef1m1fHUXtKdAMTJ3H/xLX
hAZ+glMnMCq/L1fe/hZHqsLO1XuMUf3e55p/X1fJn8eIkRn9l+KinXwe8//fRmfi
9DCrhMLb5D/DRZkQibCH3axP41N+gQi4I5nXK0/bJpWj9xVKcWFKhEBJJFV/APvd
GJmbp9gQ4ZJdLddTGem5+a35ZXi81GMs97jIxxE2nwBmekUFNAamSMVBG+Xdl5Lj
m9xOj0T5JAvmsZXBs6JiCCmg5goMB8EDPBEPaFPpCwApFPCoSzTK5shB1XnQe5S1
5huaaL2srSM8dd+ci1RM1ocgKsKOPFwmb3ENudA9vw7EFkrVMr6/UUnt32o+INxx
6yCwjdYA5DAlDnmvce1Zw3K4n0q71So1xWldBtJ0tL9tS0tFhsRYRCvFvfUDHcEC
r4U+u9ZhjztIchgzb7UWjNSvi1bz6pM1AIjbnUBvHBkBGknvQKp+68b1uS2MiPuv
Kqn3IyAhbp5d18j6IBAJoXXriKhS9ah9adD/rMrh7ioUkbLOvDMadYaF+mMNNKtB
6SkAoGRbodfOrVLBnvjaasIm8EUaH3+V5KbitYJraJya0B4K9HvPwE+Zayol/6PL
kbBVHB+GYNV+jYUzEGSFfAZVQSpys6HMLqJ8TxIn9FbHWwrwG6x/KdZw/eOEpbGV
PfdQVRY3hrwQDVKuTSlKTgVKjDFgGzijWh1pYJp+OTcFCOD1pLAQIkEYDk1m/QH/
9RVzZ9b3Dfg7Qs3EI/CNP5Wo+lJfv/KL9Qn9jhGEBXAvoZxCnmphmQXotaFFzx3h
i2qu5xd1nB2B2eh2FIuPfj3+c/pvfGK9510NETlAPOWoILh8mzMjBcZKROizqERY
mdxhFQIisUClJrtejmX0EmlzpLPK23PW8kzXi7xPhoUaxIA05f1BqWcYPr1ikaiV
TThUEty7wmjp8+1SlTI2MCyTwRiZPwHWvL8FGQ5pT3sX8VmyIyLgMcZVahzuzZjy
IiPrrce9+rjGWB+JXqiwjaX6e+ft4IMD49S9w10un+SC5PJMyaTzNh/xfWxX49L3
jn5Mpy1A8sYd7uZ3dfvcsdmX/dP/O4eN3y+wuOHO74EmZsVl9ZU9uETaoeyj71NU
p4qeCfomeR946a+vkt2UX76iryhe8rLb4PGlYS/cayDMOFdXBE56VkFxEKkdfXAL
zFgnlaBTDzCXAzUMkyjvhSFULoO4dp0y+/7tM6ccAKhUQ+lJ8/aG8vtwn1r4VexP
VjCwM9hPWWTuR8ouP+NbZKBN3pkpF4DtsDn7qy2xQjoSNSRq2lgyKTGt0u64ql8x
rQbb3fBIzwKyukaowxWclVQTdG0sAtXJb96lYvMap8YHQ163Ks4n3pGQi220wknq
5FLN+Nqfo8yrlsCA9JCgKVWqalEPonvZXFOxHSbqDztaUmQ/HWopl+4So3ANnf0C
8d306H6mMjbCLe9LatJFCgGScPAQ6C1HgoCzSSIexcciXT0uNHaEEZDKUDRVmEyh
LmY63oheqNGaRI7KZpcQ/QUA2uAaf27wAuxkomwX2v0jN8P/kqKXkB+U6bUcw8kA
GqQw62s/SA0Oxk5XEeXk4uhjZ26V7xdCssYRkKsuIkvM17OQ3LoSHUALxnz5e8nC
3Cavckz4OKdH7NFiJPUo/BshF/irt7Mti3xWa/bxcHIHl9eyoP4G6fk3EKAijRzj
x/ihyMyUSv2NItSW9KZj2yGBptYcaoVbBLY57guCILSsF3s4Uo+kInS1us7kbSWs
HBQhd4VXK1padTx90kUqferVLKR/9IAJfTnA7Zjh2+4IzbpH5V3P07cfXDR84dp+
00NVuPMCJcVDDwl+8sBzhKxA2HpE1LsPtV02sz8w3w2XBah2FWdokQW8rUj9oRFl
HG78XJYD6olseHgXTirjpqgmNiQecERPz8026hgsDNQNQxR0krMQv95cAKsvBKKQ
o8OCMAw+c+Mq4KhXc77gOiD/NUeWuoR4f/J3oWC0iBCD5gJ0J8UylF2toc5Bhfa8
TihSiB2M7NTsGO3Zg1vzw4JVN77pauvuaYgfRX5+2y2bPOLEGBgMNCqpRrQRsaWl
C9BuwSJRVP+hrW40Tn8L4ojg6zuHp0SXZU+RciO1SaRj6Ng3je8hrhz47uQDNp8I
btXegA0WzlNhJGel26AjrKBnRvMh2Y7Alb0ogVt81Tv7sE/psS70p8ulJq/pA9il
LL1w6KSRRXUVAJCKGV5cA18U2i6H0YJvM07OI+bpluo1uayKgPRLjVlkM3/AEPg2
1WYXiCKF+BhP+10vzNEj+U7ZOxQssZZLry+HyrPcqbdU/RoPmMSWZMX4Eo3P4hsR
LRcEd+FHqaWjbxrmIqFCqI4IRzL20Si4VIK/oUPeCCQVW5Q3SS+9ZSrtkxLVrPEx
1aEPR3GOeL4Zo3ujlThu9M375WuuVthnM4w0Jm7NaKyY1ZvN0lNuHHLFlZ8TuUJH
OumhPAHvakTq8pJJp4w7A7z2/mDdQQww0umMjJwBRq/rF2G2DC+4JzipeolCTeFN
wG0AADrM8HHKUWxpx8DRG87VP/dDp2BViBdOD3nnzLPgSgPc6NlKm1rgRFc1yNhG
nHD5sj/MF3uInSee3h1Zbg6lTE7OXkV0+74uzqABHVLZNYkYyC0mD9WXEg4y0pth
x7fuUhediq/qkFptn9FO6vk+3ppzD/XXMzUGZDFAIK1/u+BQru36xr6Vfo8dHnah
Qs5egfHlQZiGRuyK4vZ4I160uqLlDGReVntDLRg4sN9hWFVqZrXb/T2bjFajdI4y
VeBMHUjvaLR8Wv/OWQR0abSr4G0oInXoGQGWzZs0P3TxggOfX3Q8PhXCRwTa51yB
CIqvxjAGNuZHzKpx7djPYLNoeCND5HP3PEobhTuzuxJtj1ToiXmhs3tTnK6pV7pK
+0o8Fp0wLqSWvQY+Af9905eV1RAuX1QFq/DNlYYq1nT9lswaOaBY3DFRQQ+Kv9Z5
tqM9UbzoMtI2Y0h71fw66rqIW7BmXQ0cUtoEYyXJsIRzF8IWkaUiOOqHlCV5b+We
psqhuz2hTX7IjitHRLctbhmxbEQvVxycxx8Hva2dSV92ot+jPYLdMmo2SLM6tNtq
YEfmI6fgiVu868JlyvxA/bUSzDHPUGGYWCwtonGoVEgLVVPRmHccYwKHNXNsQsgx
mPxh+djHZPOqvxjh+NxzTal4859Bsc+2THsFlHYhWtn2Xc0tiCqWMMMWSam7BQEG
K1ZTamaT1jPIUQYSJDSXYnDFurHHiNhSDhe1UGUH1nmAeoxzSgTBPB2pvtmzevuZ
V8Htgp1yopdRF40whpssXgyS5CUCZAXYRxupv9uvE5HxN09KiMGpxwPbzVDhFYV2
IfQ1kMq04avPaCVW8rte9QXLTiyt4ofTMa8ZAGKFE6PnNoOOV63Q2IQFcMMpUcf6
djk3V74QEztozt/AkCmhi6xv3cAmK0ff6Dg9gx2N/OyIQFNc/r948deD1CTglEvo
h7cBx/RtWi2LMSDWddNaR//spUAHxJEz2cLAjF91UAlXCBLESo6vMmEZGt0d5wR1
boOy2O5rW9dY2Mb8s3AyseFHw1H92eve+C2dLDxc4SLvbHn4zAyRqUFWh4u50dIs
UvzgMfqf3qkE0s9G2CaJ8wjxxURtYgnPioRTUdnAVtmynCxJcClw9q4uPF4qg5V8
QoXW7p4P+oVGVrba1HBrjiLK3Q/tvY8yOZh+ocA4kLGxXbRdqqMOct4TGrkdP4Vo
oXtWo1TdaVgvAQFdM3kD0Ok6+9ObY4hsjlAcqI1tBqUWvw0izrAjPnrwbmht9YR5
mBfuiRqsLxdkW+KlX4+oHX+4keO3cmvxOsvOVvilbdnvzIhip/3pOi9PudnJ98u+
brPOBIFr+JyqXuAYr66Sixe0wwGcUy3f3zh8o8B5bcDVKy1I1/LUSnm/F0Ast2TI
tJIe0Q4ab4VvLSg9XZjsrdG4mGl9bXVjHFJQmFZaHHC3EFArtv1y4A/yO0z2pG/n
WZYvLB6tTVkvBl0V2RlQ9RVkEAAiouL6CKB5Uv6F127gBsk74gZ2szyD/sPd/EwB
0LWChcJOv72dusDc2MN8mr5mERZK1FBmv7JsB6gHjPUbmrG1GFua4t8guTM8lE6+
s2hnYdbqEt8+i56a7898+k7F/ku2p6ec7PtRq0xWOGNPteZjmygiwR171EThzU1A
JzdU4cIxwgGMYn0/ROYjH+Rc//70e5a0ZZa8X0XtrkmmLPf/vL1Wzt0eFzTyFJCT
uPS9hHIxOYJAPTOGIu2ItVzxVwdx6tGBvl4dwqncjkrzqCSRFalJx6tCeWm2VrUl
+8KJSos7igrRv8zuvFRTApvTSlwlte8catLSrko28JCTaqTS+e604909LorgQZ4A
Yv0o+LOHtRWkQ2ZUOv/UTkuPRIAtH7sENddLsEXp7CybIXVpF4nMzh1ssCEgQyXd
3iUcYVZR1SW1bHsAIBtrzfxpclZVWnf7XtNyIYx9JwUX2T37RbJBtVoWIn4m51Bb
7fDQsdk/Bah/V/7cOfeg+A/Wf5feI3NgIQjZWLYWBDpk/KukSwCAi2pyq4c1CItO
mgh5RK7TH5k/jmcG1rOJxtv06snv/lxXX7Z5WAA/zCvXm+c46hPvFscUvyrswJk1
JeDZAcFWSN6PTIwWMFu18smjbaIo2b7XGqDsO42xPhUlncSue8zcenJDjysfpHAf
yr/s0FS6h2KAzIZGPdUOBBVTZACZaHaNJaawIcyFeHrpNeSy2GSjSNd3fhHgu0Vf
LHLLZ2YQ/4PyZY6qSy/YOKDzQrELARIJflsRmciGuIerJbHphtSkRP7uYYy5NX3d
GGa5I9xRpAYXpvqVWS7HCqsCYULam1pDWWOvwj+uMHKOMhpDOGSdUO4j8FIm5IGO
yMMurH9H74yxSxairhNxqe+DvXwcC2g1OX9sjfHrJy7T0lEhkiApiJnzMmRSY+t4
LmUGi+T2YHVqnMFFkAoLituHr8dpdYeXUOppH2qIZjRXIrBjhtHEpdfqIlfIy23K
U4meI7ZF7zxMXUBRIYsnXGnFk19ni1Cnm131/t6kHeDBteDcXXSy/AKW/tFKI+Gv
M0GJKC5+RWjh1IM1iz8aCRjySMp8G4cVctTkGmGmE68ha5Cc7v6glGWiMyWQfWvA
byucDTG8/l05IxbeLCkXjQqjG5hI84WyAZ1CFvEpYE8443V5/m3qViIekN9UhuFe
Jh2hx0ZEzxfV/6w9nC3EIDKForWPZK8+Ad7x6hjh0kvvoNvNTjjQw9JMuxRyZ+b2
TzbWjTrRN6DoULAj8RAFBBhpdjX9z7O2dHbjJQdpy0RqsmjSpTcUMO73PZz0gGES
QTz7/jw4CU2J1qTBpkav73lm4Me1iXiPvna+V+4+9iGPE2SEp8xilYgj5W0/8rcn
g0EyIox1PF1rL4VpasrncpUTkh2FZStOhIBbVLo2ansNEZS+Dg/SP0RMlrmSMOfM
Qnrjm8Ki3zbwt+MUqM+NOy1tFe18JDKmgH1XM9gcPRiXHmKgW6BLciD6lANwMMXx
cN/XFDLgnyhaJIFic4xOQqyneFqF9bq3honeaTwFNLn4QSqQlBdXIuC7UlyRgEgc
jzd55B5S9/lCnoX5oS0Vmtn1u0gLfkhbjVI0lniK7CbEkdwh6cl4qCXOqbe1aQGN
tZydvmicqxPihMmm2RXyIK8vvj0I1fdbUesws40dfcFXJfHOagLdYEZh2PNr/eHC
WGsc1qJSK8Mk8fIdxLTKbDwhA6B+emaPZXIV79NVmKYJtlJFNm2VZLc6tUAG0YNC
VO4S9HZIVsNSBl7rjwvL1h+6bjJdMYKngFkQL7IsdgbKclHOvtaKrTKUEN+nbLwv
t9h1HXKsHdS/k29c4oFW1pSkb6Twki9OJk0h1DzyD3j5TrdvOZr7Gq9GrBwrtvPk
2Pvgut9C6O/QZ9CRoo+tpYIt/NLuE/JRunEwTrnZLrubx8OnfMhkec7+YdXXQpdv
BSs3Q916WTxSCF1dK5XiY7j2f/sSsF/mO+yctvEuazpPbIYpYDuyzXrrlXm7JYtg
3GlMHJy7FWnMime5ydtEBDtJ55HjwUlFhVdnKZ3F7P84LuNGcHfdq4GS93mXouBP
75/E7+Qt1ROJEVqn+CF12reaK5JzmkxYKGsH+3fKo3GFMUvKN5xXVpH+wUJEN2P7
zquGsk3umgX9kARIjOj5tcreK57tsmkyRigpUSpj1W+DbHqmUf+EWuXwQPkQRWzA
sgJppe44+eGgfSvLU/oK7NQXMY7RZU9+T1GuJVTEOgqnZVlJuRqYKJHGrH1enZHk
36t3BYpRkTdQMIZIDPDfHQavsFF/ZfUGCBMcjUueyQdIju8JmMhY7uanMlR4bFAZ
PwvI7vdGY1yI71fdhisDm8a1ThLPghvbVa/XtBLkCnSlEUIDLbJwOG5one6a/LAW
evPeGjrdoxJ611WCOvqSDrQCHxnkBFr4gCdGYaoBuHdcx7sgphC/PIfGbSHHEo//
AnlTYrlGpt5oq5IEer81emwmI3dK27eidsP5VfLUX6uGmL2p2MuY4JX87ACtR1AV
0hCqAd5LQ2Dg7eAj+mRAuCLvO8SWmwgi3YQic5i6Z/yVxjhiX3I2M+xMQm+NWqdF
IfnHll8O7uXThPMZiEJ/OuMHSs0ETKpRXsktcxhAntZ9FXRAHMWyy+qHOgB3lO1i
d/0tAZixeiXI7YRJOkHrwNlNd7AHeAPNGTP763dfUBFoP4Fh1m2at8ml3FLhJBGL
BpvgZiRAAZLtA0Lhgt2HCZmWRkP7IupBxZXePRqMuILs6GTvQPPvFOMX5jQFCeto
WMUQ2fnW7IV39nrUISVN3Ebase6GWxsAYNlJIiuvXlmUiq3VYqkKi9GoOhA9Sf+4
kQ1jmSKuxLvnXnTEc8p/NQl8zJq7GrVS9ymwBCZe1IRXRPYPgh+tB1OG0HoIURGp
LA9whfemjU2DtaLXw8kRyyrHFQY/YpwVYhwVOkDnf/CXztGJGJWzNYYEQcZhVVw0
WJjbIYbbKmOdFy+n0VoCRFOWT/q5w+eBpYVReWISljIsB7kVK24RHGfrZC4Itc/j
ABlwEQBgkRJoQb7Eon7//t1YgwxFdqEw8i1XTk3oN5ml2J6yidlUzpIfHtj7/cuz
UJdAVpiOI4gduI5/oU5DUdkzmetGSFV2PnI3IkMQPODU4+r4pLIaIa2N04oKcwMA
uNQtro/Uv7WObgpkZ/Pkg6n+q7MfwA5HbEYO1pBuSizs+EhVMKVAYyDf6JWcQ+iz
wttOfFleFtLwVPil++d9S0jiS7M92o1Nrx1UiTIcefp35l96KNMK6F+svCHCFUBV
QMfQakH4cDOZheWWi3LlpXokhZkNu49fQpPdWBzo6Dc9zlhoZ8Ip5jZ57maKg7JB
7uU2jNy/6j5B/f0v6xFb+TsSN4A5ga45+lyErGG0d2NzQih6F+Eej2RZ3QgjClmh
6px9g4HGAGUS8KWm81dm2YNifIiqytjxIOt1RB/OOw+dKfxvQqxU2NMyvZTIWEtj
lka0qlOY+AmryUfxF7YZo6+9RRJGV1hncQ7CXTqJqGX97tzX0zVO0x69Wig/Hmrk
0J2Ckq8aiqhMDTLenU7wi10WifOnNxF29W2/r0cbMdWrtkdgB9tGT5RckTnmorkt
kZqRvRA+sh7cS/IHy83SV69bsezUxl99GlzYVoD6NKuquL65euBLgOETlzr98h9Z
jp0A7r1vjZ3hX5qPgzekWZ5M/yaVWJKhAm1b2vaoA7t6BMJGkx95O7WwjhkwFFRZ
k0W4sajN5Fuf9YiyuJpiHYS7fPoJB6r1ECSQmPckogAluqwggrMfakQ8BMd2QXnv
6JaimFThAEgjlMl5xXVEAoYY+R6bSbkdV45ydMNIgxzIoCulTJ3dXaJanH0fVXF/
Xsz4H6bwAAscyprFuXUVkoOUKOdbxC/E6RMldC21XcvIW4SpSzA1XnIudNKYKj5B
X16Irup+UAonlCvewP0L2kAZ+o8UfrJ3vrc4wt47quJb2fMLh7PfcIS8jQMDXVZe
i6q326YUEi9wR/OFlql1SHQh+b5MugQvcwelCh52GrA9W/S3j+aiHMLcEgqJvdj3
xzeuITJ9oqwYJicOVS1WP0QlrNaqaOW9Ked9fRROauOJ73UX1gPuuAsjBfEgc3zP
LxgWVBk6sRKLfojuqBMBfjWpD1HqI2T89kL4OZ6phTV/dLEfPlyuCpy0st2v9/qm
7ONIPzDE5nsctvg/MFqflJDJlJGmuwZ195/oKkmXnae6INEunw8/Vyz/lWgc+6Ao
9YfqZIZ2ZFddJ44MDhhHwZdtNSbzpS/CQcp3KyFB50Sxj1EyFRMPn53490PkQ+Yi
t+lYLbPhG6T42KpWU+YMSRI3lJsi5CDVcroWiwVfBQofYvdiVziNWC0sDw3OTJx2
ujjuNxvjNvenB9NVNX9Xz9610SV62ORl9ytV00GJoP+oQQTAJvYO7KR66zyoyVby
HdIvCqJIn1XLpyj0epvotsoiqJ+x4vKl//i2NknVnbtyY/ISnMct/s5j+iufrsiv
mxTzVmP2ZJjTS8QWXNqMUzvlWNhJfXYWLHO/zfUaS7WJ3plPs3ihjjsJdLRts2ML
G4M3L42lIMfYL/HlU4RLgNsvP8A+KZ21DXz7swf/ZX544TQtfYcrEuYdWtvZVjeX
3FgQU5cbX8iS29E41mclH9i/8WrL67uT+Ykt91FRCBgXgj32ajHECZlN2TS6IREb
StLEmashDHH/KG8xPCETooBED5QdTQKUB7hSs0dsMVyKPPZZMYEtt12lvV8KR6pI
m0Rd8RbWfpqdVpkYuhzgts4Vceq69bGtZ5SSwAucmzYewr8bKONvDsAPTUrtBFgX
X1jz95sJJM1TFOadsAS7a46nPl87d3w592il7a6q9kS5GCK43EuijC74N6X8tXOb
z5yQknz8//HjTgTm9jw5/FfCfaqjwx8XICK2/FfY3RCUDrAmqu4FE8aMSXb8611x
E1sXe8gz9HP2x4ghCQ64LIOCumqK9VwwEcvuznkTl65uWZUcEltWsIkEz4Kvq6bx
90FzLZH1b4A3ry3+ng4HqfWzz/NHK6XH5yJMXDkIk+hGNIF5u7DiNyIODuUs+PsV
/Drb/kNnkx1WtaM2hdD2MCrCFxLw4xT/zJs6hanbrVQ5ImA7bX/agNy447KNhld/
cuG9v06FpKXhSAot7ikArDR/GpBYNTqQLNJfoOFexnP0XmTdMe+H7q/l8SDie9Fw
JIdbb/t7kjVQvozvMe6OSVC37zhu0ORRHNvHZlTnsrk/JwOfD3/v3YVO2lvt7a+i
CamnSnhHkSuAi7BhO1fwUEbMURftCYz1hIlNNKOT4tvzxnPQSCLx0TOnQYnY1SNI
KXrO7W3VhvjwH2UVS1KZ+9kFzvIqQg4hgVtaJcqD6dlej1W2XMW2Jua2bwuvb0H/
27a8+kxSj86j2aEG5p4cq9hdQ0Eyv8RKw5D/thZWO6H3jHakL/Y/CQwFCEukGarP
TlKi6mhx9UGfmQFLDKDAYTX+KAraJKD1GLopnqwUU1I0/pTvUkm6sN+rB9RNlT15
UcQIdm4NAfykARX0Nq4B+pBbe0fxwmhzqw2x1O5J++LztMfadoSxHHr4hXnJUXgE
JYi18kUpO6B4i+Zwj8f87qHmLll1ZhG+VEPNf0HwRi9RBYZabEVbxFqnjMFGwlk1
qTiXO+TdY3eiezPQbaBgvJYc2f51ySlzh8GeTidmKPptcWskC3iThsjlSbHDHA5H
5iv7+mUoeMAYQROCkYPExgNINkLVRze4HnFy08OYgK6zzDyDM6NXMWyEIFTlgYFf
5IVKWu2J/cAeIGOgh2+jcZDrvdTKvjK7VGbT+ZWbt9rc2TiB/eyhZxNjdWVy9AEd
LnXmJe0rIXkwWpObhKO181FO2i8JvuTO4srOJz7/gnvtNlptZ2AO0tcDQkKgT7vc
VEJzBkJMmUOr2zes3iSIYuMhfnGCCSW6QFdB9qeh73176XLQA4TMR2iz+G+X+CpB
XcN/FlBo4EDp9Zlt4Vy5ZumpD1y1WKEArW+buKXooi38hQXkJl9OEZKXnyL07h0F
9DjRNBis/HzCMOxFoYJzbduVZo338raF7ZHZO31wWA4wRWVbxA4WfU8vr/bJ4BFn
R/Z9bq7lrTuxo5wdZmHF6KmN2qaaxN+rj2j8KPpElQ6qFZBhy7xRaaCG+i5E2NL2
TI0NAPI8rWajqUZCOMqyTp1BSIHD8WuHnE/sReSgI16ec/4MGHWxRufuXqweW45f
VinKgps4AxIAXZXlmMbG5NfvBzM9oIbd+hJQsZH9JM4YJn3F9o69TaM5MWad3ogI
pt+A574EdDQm6zjBF09lPTMAqSU8SQPyF4PH2l1M8524C7W793+hL0djBi8VyTWg
f2dKEr8I5uFUlrUl5uzIzmHEzLDEQh4fyz/y4XKKMfqTtwQKDKXFtZdU25nodmAg
makeR0OpuZTbH8oe2o0TYFWBBKgVPklcGn+4wrNLMIgMan7lw7nsp/7o2tt0EwYg
t2fKsVRB9oCQeepNnCAJp6QCtPMWpxF+KaXU8cmYu4YFwvEZVfzZkw00Oak2Y7Wh
ABgPcExIjcpNlR/1w+gkzk/2y4CPquzN4ZvcV42l7P2mex7LpOnJE28c63mye5uy
opVjvPX2BZ6wRk0Pd/EM3c3B8WGTBdkfM9EBRmUom5/TAUjPBeEhHqh1Y5T7GpMU
xCEDZWVW3sNg6LKJgEdMHdsIsV2J+PmzTTZRrHtQ3Qjxj7GAmJuA/3lY74vX4y4S
7yZ85yAHhzRq61IMHuogVmSwRrzTv4ckEk9uiphYP+Zw+XU/vne1SC/s09bDuetg
9Qtts5RLGxsvgjqRogSaqCNXxQ5FUgd2qZaTkrbUWE5ZAhLGU2UihDEsBwYIfrIk
ZG1UDw8l2pri6VZBWQF+VQVWAnKbOORdCrwSFEE/Vk9BzS1ioMnNK5CxRg5epdf3
is6EskiIFbU2ITgnMQ+jZnwmO6RiM61+iOAj73dkhPl/lkz6v0z1rVdW9ZIg7Ixh
BfhWdGy2FIMbMs6uzEkUSZMwB/xVvznkRK7gWDNNjyakIyTg4QF9mf6mg7Jza3/0
7QNM5V5+Qidv9v+iFsb6KFVSpFe4CcotFvFC1jU+sDWXMDSijPn9L8U9MQaWwzDu
kZfw7z+RprU2pTfPae5DNHqOYptK/g74cW4zJqtJDJpmAEmm4yiKlOZ4WOV6yVVH
n/UDT1HdgVG9c4XFyoLfJD5QQLRFUC1XMI6fYD43xvRfg764A3/JnYVuuMGY4HMm
rvorBENeFCGEiTcLF1R0k2nwwkQdVh9rygQTtRnQuKnN7VXtOKyjOvYEWGXS3RHf
SzT1rFDhOkK2JnuBXfzBV9UsgJU48novqXptb4CZ+OVgI3vlaUglrfWueTUheWvt
GE29rks3tF8p2QA6OQ3gxqgKwufu2cgBo41YNHUqjhZdhwqMI1icCzxCRSzio6BO
oR8ttlJGYds07eWntl/BhR0UIMwC1602L7bHGTYXDPqaX9DdckUiYa+0F8ui+XDO
PkKyqwTrtvaBPoxR+sPXgZISxYaPZSkxXQm390bX21OzjPVVhRo5Md6z9BdPHlFl
v3C9lQR9mrGJlsiQtxZGyRzgBkZ2pAhDw/U8N9SBQ2L/TYehpvSY0fb2j++Z1UJy
xV/5GvK3+W/mFIWEX0ZFcurtJD13tZA14m8zvYokyueh6QMpel6aG+HVk8vbsDPg
UjyW1gPhoThkhICPTobb4qqouPVo7PhX5DkuEf7sgfMuGhJhhTkccL8hVqsfRSvh
FWoT4+mHrOiG2VIujKHCZ6iE8kNIIFX0McJ8dY5uJomAKsvXjieN7YQEgApmJiLG
acidOCVHPqW3npc16IGtmcinvLFVERFytJEjQ9kgCUvyKhnW/LFU5LURyJ+Y7nkk
rl7+fUoP2SdlTPQlUAcRx0h1EQfthE2Lf+FGvAL7yIEom2Ld4Mnuv2qlo05NEMF5
6DwCsPd+5r1N1FtINl2LOWBXTvrrhxelrSziy112dH62D+jxSzlU1wgPWRyXGuro
SZAZK2o7poakWKqaT7dbJisGmLOeHKEpkgyGWhITpXDFo1SBm/EZJt0Ty/e21P/4
K9TnEhnpE7JoHg3nOzKzQajsyN5641Nn+LLMjvg0ov+l41zwWwtb4EagCTt/KVUI
2gcQnsupTQRzBG3P3ZnViSXFaSAsrCjZ8lm4sb6djUJ/Vl3UcoyIK1VtjOiGbWii
me9fdVHcR5wGYWHHrBCnA0UzPjUKxTqpRLkH6+8DdxVt9SG4JaR89Je0z+QzhV+m
8P8IhsP9hLBluMma7W7HK2Cfj/CIeCaZuvTS9H1gWHAlEqB4ao7/HI4wGCkGlhtn
g8msgGdytGLFkGy0hfFhuLEbAWgHfQdTipqtywTfw8EVHYO61FlWPbFFElWb0ygy
Smmi9LQWk+0+zsHeGOc1iLdGf8ESW3ms5GyJWmDF1nIdhsBUM6vHYtIxNCB4DW7J
CGeNytOC6fftHBc1y/o7iCnJw1Z6J0jCutJR3sPHCguIH8T9T3zHWFlMaUGOcfuF
796IzO/CwplIjdtMnFJVBITfau2ANd+vCgqYu8sh+HVUAW+hJX3WYcL3/S2ojUFI
bjlw2Itp47XFjEDXJ8sEYcKz4QiQOD9OGkLhSlzIsW7xmqnVQTvmLwMl2pzA3AsJ
qJ/XSBKSZwyRZlFDb4qppY2MZqiRo5gY1yHCTz+1t1y9grl+aUl9y90OUOL1EHbh
c+lfxLiGHGLBkBBvhI2fWZRePa3+N6RdjP0tPhh9Rqnob2XJ49J7j3aEFiHHj6d9
QgzyzdjYrhypByt4F7fY1KCl9aQZC3Yqr/OE/ymO4nWY+xPIoRfw34+jS0oTGvf8
5jy3ZaaCJoGmAMWtSFbMl+nsIahkPEi78L7iFluzNjeIBOBR+L3WPyjblPQ1VccT
SAIU0izG63duXUOj/HHrOh9aSPniI/tzdjPhBFncBPJrxKbgooCnmvuoEj3nqZNs
lPGZmfxlfgI8yUWLWhRS3Xm9b5gg6k2VR6vUAuEaz0IrwCo0UroVh7zC4yEHDTj2
xbrIG83udlRE3tsAdisD9CuVMh2Txc9GlKvp1c67uhusc1YT90J9B7xa5P1t4iwV
30jNyu9DwswPbizHIcuS2WRnjjiW3o6YpEhK7H8W7tsr3cZ+AapfPahgufWW72u9
WlqXJiSpHh0bYJ4LA5gqhpDOqYIBWIfJKDlNQKXQJZPyO8hBXdyc9uLOSuZMHCPS
MoZ4B5/lj0uQbdCpsobP6dBrcQypnJmQJHodI35acQBfRnQRMnFlrZG5abnvkt1z
zDlkiCB8mLnRO7GkecaM5in1wZ4Wa5aA8kyNniBcfd7k3YjA3SdELNtFvVp0nQ3Y
MnP+hyOr8o+loxcwQJj0dvWkgnTiUXWtlrVI8ZlLjooa7K31Y25XuA17j5Sc4NuY
/lXYjmJbw28ksHvvihTVmG3A23qK6x2DqZ32J7NJzU0gTLzGvrncnaCbtg9B5o9F
nOoR4FxQyN+k4owv8j58T8c9/KPfQI5lwZxdNHL4qxSCsgMVogd9KIYIZ8F+xghb
iTRv+kdrjXvAC1Yb0JSJYgOdGZtxjj/0iG+5Zoxk64NGfquToTxNeNfVK0jdMYpC
mQG50xIs4KfZ4szFJccOeTmqsbkFg7hhf0BhcN5nyfYM382zFMc4wNo9D0eJl5hJ
bTPOjjZhNlcuFykQ87xtO4SrrqH1Lpxr4sbP9POVL2Nxpj2pmi4JakPMqx0JbOkI
KuRuwP+gbW4GaANUUlvywyxLR5hmJ/dbP9xcxfZH+2rv7KJRFgdIgf4YAsfz9W6z
vghlS1FRfqWO096s+s8yUGQwNx1boCxC1Jqj8/GK3DrGJBUinNDLw0jTXzwhho31
Ypj8tdZ2/AcbgEJK0kAt7eniT6cuHdInLmSLiIAvjVE/iGEThf9ZDF3uPOOJhuTF
15s9L7LWm2oE00azF9c896pVlvDQSLvqkT0Y5o7+MKGeqQdppgxLGcXhEK1iJBGa
3iOp9/6lsQp5VWod5vmYZDw1cA46jhh5Gy0caOCTi0hTign855ZOjB/Rq2gJ5PoX
olVhQwZIHvaSd5jCSi6+MypqR9B/7VwervoWTwy25uA5ZK4lKNiWXVOXuglYIKer
Msge/cn9btToPfyFKZXsGUEAKwNUDvGcpOp8nY3MpK8DzE6X3Y5kU/hwW6+Yuazy
I3mezv229W+nuYF1L6jFv425tuAfk8B3l0VMHi6hFXmazQgBO4uSUaDGlK55eCxY
eIFJGT0lb6FBpfVuwN6aBR+Pv6z3vXL29ztbUzKGS2HtZeoiStB26ZCEwg4w5evN
0Y1FekP/6tCypXUiMoj9OrvD+vW6i6NWN7KUuix+Ppeh9Tv3c7UiGN620qSdzyHb
L0rJ0UCZ7Imp1j3j1Xlr1B3VrAnsYO55IgN1TXA4SZERWIgEJj4O/D63qCyXYuMI
6BYRFREoUQotG+iZ65SDLpgdKMHB5IDkDZfcVr8E1l29g94oPPQL18xcw0/rk9sY
pIXoPdweFQypdvITiIGVAn2Jk1BchOdAOftjQIUeWoDs+MGPUA/ZHBTvMQ76c8WR
MOLaG14OZUN9swSQD3vmzEkcmdvQrQXFYJQuZ1QxIDyUCSfhIifdX3gXLWO4O6zS
GIx5UP3GvziwFZJynZ9rJaBNT9I5FyHnp4jjSs2yxXvZ4nEqGZtx7wr2jMnPnVBS
36rZGTZvRg9GFElAQw9g5GJoOLr3N4A4w4JC1U/S941EAIlI5JFeBL1xKZTlDH0J
Ic3tpoXDHHW3r7XxpvhENNl6KrNjGencnwpV7C2fvZuhdR0O8OOobtCYPbqeBZzh
2LR+/xiYZAvOnA0ghCrEcpoNcOVzHgw4CrqvBzXDKGwH3xxyiRkWOFPAZtmLQv/J
QygVNFNXe0UqLf5yW4p5gMI8viqWAiA/DJZG6ASjOEoYNSGcaqB6Mx0NGYmA4/GR
qe7NTzODwHDf5MbOb4OevSOerqqlWPpCWP8zGIyCL02lRFRGK/ji7ojisZJgdRUu
Hg17zMb73O6255enW/KdmcQH5GnWoYTJp1uqRJ4ENB6KLBZSDpV/XiAPQNe5nA/K
PsYLMiUkKii6eAkpiLZAHUA8XiuFMuWnBnZlth08Anhv61eECZdGIfLKQi1QnFmm
0/Xde7vF1a6O57NX/MW3rtnP3yA0z8qty07JI6T1KFEKeZPLDV2D2bpwNkfuKLAE
Q5Is2RtNsFhitGE8eqAVZjEy7kHEfHJRlSbiwFP+tLw+hoduCPNd/aodcEWGtcCs
epFGkAg2wzfdZxtfzGyExCuuAiGqhmtNSwrHjt+A4bTTvQfL1K2iSW2atFex4CfW
d7IJsyaMwTjSobHbxYqFV6ORdculHX0MwKJ7QUvC77Pwn0KFZnHSu+0bBRsm53hh
VGz8gmNPh5wKM5CdR7egs4ZwxfAXyx5F4rid1IPNgDkDnCwfJa0iAUL7HkY9YN/r
MKV0A1dmzJlHGrdktPcu9ymh0sTBwCTuuHyWPALe26RC22kVpeuBZ2/e4qf7Ln2v
wWRXoK5y1tRxG3QE7HIDfuJv+IUCOPHrfQWA5JkxvCjRH1YGirOwdAzFJS/MBc/W
XvbrzrWo3Gcf/E+qKoFNC/ilm0muurfDFEIrHHgFi1uoBnIjrNZFmt/nhkinLCSf
e4nryCI9Pt5dfcv1dBYk0zm0UgixL2mCld7HxrK7p5vLu19BxHry9juMgOuJVD+/
yDncLUCdoY/2fy/tslwO9IRn9H+66psXnju3SBjNyCH7QGNK0/r2lvMQ1071xxfQ
rMB+RU8P7iUBPbuBMbL6bC/q2U7s//Gg9Rudf2vGKSXOiJA28LGtEc3H1Vz1ln7J
0VpO+9PRJK10lR5TR2fzXsIrteBeqCSGHPjGokRohbXUeYrYflVtUs2zANQGzAhV
NTNJARl+71+ptGYkIIo5edqrdZVJoKLzJNrm3hPk16Gh8G+0NuyO0uJbhGQuOoEJ
FhZPpkFB4x1rVUgisSQi1lMzT+Bbg5SUGIlWylKytagMbdk5OIpdRJxNE/PI+msJ
0QsFjnG9Cji8em2mHDsd5oV6YseVlgfYZmh2/X+JZRYDh4LLvlwuhSGnWk4JC/Ip
a2Z0cmwMFrCQXWE2mNvqcRd/vjDSYyPw0zOXdlTqEI5F2ZKp5Ibo7A9Of+MK6QIT
ZtjKfKeC2itoiRWhcIxiX+upWkMrYLTishvtYWqzVcFySXVvecvgWnfoFopYRgHS
HH9aNMvFJ/a6WkbYqWeYcA+woyj8/osMlAMAfc/XVV3+4wgzcmO1U9P/1ka0WHAE
Fc67zlthWJs0C/IlNOY3fmH71h2ov/I3PvVBCEctKRHQhlb2FPIZOUgrK9xzye1a
Vr1Taxappf/tkRLPNDeOwPy0VBHbPckkZO7tZBydlQs+zqOWsLuKksL8ookRlnIZ
sV+5CoMW4k+sbN5OLF1tIlI73efHvtCqaOGPYZoYXC3Yvhdux2D03ABfeRbGB/lS
ww9ydplceTAu0C0v75kXoxTiUjqwJMeK4o9RrkbLGhA6BZwECxpJ/Qjg/J9jglbd
hyvd8Z0zMWMqwJ54ly5rQ9G805KhdXvCVQK+aYNPnPXFxFAA2OXgn3eMdUV11tVA
tU5/FB+ro/z+LjaApee/x/53sM09B6wUY5hdH3eYl0qXtZdwFreMO48HHxffDqll
/yhUZiMagZvTFGhnOViTDhO5vgpbVs6cQrQmrlu/ujCtwK1fUChJqnMc4VoaqI3M
78q2nQwSAJGM0RZl5tmSwUMTWT9pbOopY5MQtxGQDuNVITfS5YPGxegYcCpty2Ge
6+ianzQUtEOg6VAcjpL2DCrcZK+VmF1K9FQ2Vhrl6Lv9JIiYpE0nibMrY+aj+0Uc
DaGs1KFUp9TZnagOrdpjnJvTEZT9d8BmXOzDpwmvE7nfJLTZ1f61qCKXrp9xvHvA
w1ITOjS2cGQoJvB+6RFYn1MKke8PaUCFgHwqjiKOGGVZJUgVCuVC2iqmVSWFhess
ScUnlVY6dg69MpS/YjyX3piBWPEV4lb9vtYGqqzOp4GyfcK034vYtX+p+GZFO+Wk
4V5w8EeMo1Ld6kPdpaepFJKzsz3h2MKwXJllIuZPBThDLjvIleoeMbxwuirnBNEx
+ywHku3I5MWYPPQWoYH4IGfxs4JnvF6zfGPEI9BK9wwN0G76TXyKpjMg+U8CQKa9
2gA6IGOpAiYsxbnMvOnK/mlsCeRC9yt6AKjxqzW0cj8GmTMglBZC0XZXJHq6Hrk2
4mYV2kplzGkwFZ8tP67qjtZ9WnTGdcgXNcMDOQcp6Ks6waUarUgVM/bmEzHkzVR+
QfwFscK24cqEZCCb5+5w3sscftK0aOUKSl8slQ4LTFX1HWsrKRGMeutRUtbS6CrA
9L58LNS+son4bSjFP0qnr5I1CdvRrlWok9i/cTBWQM2nWP2oc10PokUukCg/dlYZ
/2BYv1CZ71mSLJ0wWcfAjDs/LEvpl1h1Si3xIZsURbg2sNTrtcVaA5nga0EmjdHG
Vj9IHVJa4XwnTrE5zUQ0lnCpDYnRObAafEtczsxsFZQuyiKupvz8fxTlP6/gRP/Z
odzW2btYdqzpdFrWhrgG9n0/+0AMgxR6emBc/30ELd4D/+hl2CcTP57pcglFdGCH
x/AgvTLYpqmGte9HkYUA4/FpSUXCjDKn6pSBuZreVUYLQLHFlTXTSBmEQLxI1T83
M3K4kpabAZozHXGsKJL77dll35Gmqv8g3WBzMyEyKELGlIFrrtRIge9CXn/kpkWM
gTdl1T9/f86sFMOB4LUuVCFzPK3AZ4OlvXvJauhHmja65WKnhiQjyjf9GYnRZ5af
yQ+bEL9Jnnx2n1elQulezv9PGhU1j3f9ow+IEJf3TFUVwsPL1Rxyv+SkDkSRyQp1
6W32jkMrJ2b4eDBH2Qu3n1k6wcIcCSE9SU2c74PLBfpAnUVCD3Kxl1+zKeMzpT1I
N1ZWYl3Avc3m3o1hSRjdL4mZ41hUELUFAhlyUTUxuJbE7nDSmulHtHyNHWGuxx1x
CALStns7T3zrct274w0PMgrFt8lIDwe1uNpXcDAWUVfyalv3hYkZKbaMcIWK+R5z
mRrpZGL+dWJO8ErhbzM6Q+wOCQYB0GbxzSSYB9z3X/Cfn1A56MY8ApT76vp4SQCL
f3yX3m8Bs7imrjFsWJfz/v4f+fgsAvR3/juHYpHDA++rXCu/+9xl7teuDP6pPFdg
lPA9qVoqf1aTd40JJbXzKX/CZrV12EGdOOOD4WYzadjQJyscxeUKvGVofN7rL3Uh
S3ywjwXWSvN86ySO+tQZ4eWdu3gs/46KetiXTp8hX1TTc0cNvG2YJOQ6/vKIIp4+
h9lHl26xP/n+puqRwDEcxTKLujGy3/W4CvTjzmXqNPhOW/qoXOV/g2RXgkxTs/QP
mBkk0WldSDzPfpwkUn/aZXRAKgwZ8hJCjlA29XK4Es/eGNyuBhrwlzsiLtmPb4St
3Hbup0uZPj/tXphKs+KbRQcIwFSOD3ZQVN/13fLYfjmWLPBKsM66mvMr4lzH7eY4
hlAWuDS9ipuDbTm7AY9fY7BZF2b/dSZzN2qHPmj3/btECbsjnHgIb75NGx9l/I8o
FHcbqtiHqcbCYwcjStqHTw+pdAFiVKEnKrE6XF+7EoE3o/gHSjXcQDHnKALsWYbY
mLUtv5/qiBbNrf1748aX2MMcLoWx1wuV9AyU6ZlZbVZGO40L1dTs39koEc/xjoHz
m7uD6jBGxp83Ay2ogw1ovDNxgS0OQkZkj9Td6+I6viz570io70B9Dvp4A7ygCAA9
2ddNpe1x/bwNPWg78wHowhYb3V29BD1DZpvh/98vPJvTKzLjBu/m5jgTHskZAcQV
dlGDDS9XJrG9WyBX1TkjlsysoR3tpRSpjhdkQUO3kXivI8326QRo6atwpcZpiytK
zTG298x08oU2y27ZymwO3crMGSjn3fIuGXGo6os8QvhQzRgKamBBhzH2LhUffD8z
h/XEPP7C3AAZyAOOSxhKZEf0VQucMTyxDok5EL9eqlGUuJiQ3qaAnq4MmL8fFIVN
ao76UcccImk8bx+w7uYYk4GHzvT4RokqJnOsnq1CeGyV6/lyik9TW8Xn7n4AjjPK
0rC202us0cm5vTK0kklwtWmJM+Sxk5SqDpPFG8PyNT7Z/UzxNqi3SzZ0hYJwQD92
TAAuacYmJUM2t9ryiyGAomQ2lB1HMCU3hTfPkNVGBl8qzKJeKzzIrxIxU1G1IyYq
+GIccUxABWq1SQoWl/QlLkdptGUUmVmlVH0bpRIwxvrfV0zo46CBc/NSi76K4wvv
fxDYUk0WEdKce4u1U4b2gmxdXemMx5QyEi0fixFa3eaHKqyslAfsl2XDK07iemsS
J1orfllS3JrDau+YqHB7FqF3qU64N8fCPEAdzlfCWJBwV4sBxu6mV+R+xD7D/VGp
87o3Ka5djqUq8I+A22/rWm5Nx0wlMS95H1TYhQ7gHI5A7OGjGbdI+kUBTnVw3d2i
GVr8PnsAl7vCaO1Cr+zvRpbTyxFxusTz67JaIFAmJ6ZM0B74gy1gzj5VqvYMyGpb
8T1/99pii6YfZXLyhHOGplbHyWph6/idFk4JodiD3A4jWoKrl61TALF8Nqf8s+qx
JaPuTf00jPsFQWcv16HrWMpgHpc4lnUwJ52KoQUxnnmBBPhznRtfa0DIWzLpHxfv
PDeLbQ667j5ElLmuIq7o6FsD/4DqFCKNzfIR8GRSH6T5hb8OklDptlRqc3hj37ak
wIYqdAKULMG5ztgn0RMGEUxyywVlb/RM7UxgHiOmqDck+c3dbku3SX6ugl0/w3ZC
KaTZdAecPjADuXvsk/c49nUA2h1+HyxgcyNN4SmExOC/9e+GAx+f/iLPnlqpuwDo
iWXtuzxGCwLen64NMbyZm7leklE5qm8WWSnv7C7smm/LUAfJKFeNvZIeHki/vVNt
xjbGLVwjLyNnJuLOaTiDlJfdicwSowxQS0aSKNYM+7CDs4yKsl2H0QM9gvxh2k3p
I2DistOUhvud/PPX2KqJfcXL9a7DLA7wlca8/DPHS/3AYNSd7Po/JxTI5QlGVh89
FUEfsR3MuXrKkmyHG0aJxA+453y14qKnA1BQocunRSuN3Xm5npm8cxqX53MNaBHN
SzxGffYj2Hut1imyengG7cJ8/6KAJkXyjVFmIVUCcPZ6hoS/VMDcZb6uTq3OK1N3
W1xM1qWZt5569Gph7fAWh13CNkp/c+IHRnV9kp1dk7YpLayLfpt7wy0zGc2Bypei
9KuRpw8uHNy4Bmct3zf4qaNiSwBS/zvGMYVZL+2YFAatmUmn6xunS+VF6C7fx6u/
6iG5/tV4i5pFZmNwu6yRPlxwxncAlllhI01bIIXpSt1PJCOnFnVL6x5ZS6iDxfKQ
21wEyqRKbYgGtZ9eRYqbbHR7MkHFx+fXiONnZF2WhAN/JZqPc/zH+hvlQSNST51I
sYT+lCQt2sksNo4fd0QTsTSkHxfBxgydmFvglxMzESpRTW2qOb5NkUHiyLgc+Usx
GN3dQJJSrqVTb58pYSwAywr4HdjcZOo75QIg116IRrzxEgm0TFL1J+5dJn7gLwIN
nZjMr9uCKEGjHPzu+dyVrmzhF1tHR62V0ICwybZdyTRk44phVfy4CS4f7a3bqh+U
SF3aGfRYVGQdLVuVJmOCDF8HMMiTYs0MN7ZV6dyOkFxhpYOIUQD8YQaDkFPMJugs
DnedhalKD7m+FCIWDCYY/TUbcC9VjtNd0U0pKgm2Y5V3uVjyAEZkTXS4P/GmKyiT
lBZ48mZ9h7NoK/Jjt/Zg/AM3io6YTwkKqg6E/2MvkFvyBrMRWE9YYTl+A0I9VeA1
823nxYP0Yz5a4c7NZMg8ouh5/7ydtfI5K43e+Dry6qrYDwT52qQ8s2145U7I4u7v
eQXjeLw78uSEsdc4CJ4HbgLgX/YiFaz12aw0wNvdPDhMSCSyTXLahnQq4m5Kg06E
BaGFglSZGm24u5vr8H8U6udYLakV7JXUGRD1I9LNyt/j8j3oQNuocbg7fZGK75gQ
0xWSqrcVBhiLoNqwPidFWGTVAeNFpKdsS/k8ijfiWoQYBXhtb30f0j2ByV6R+cxE
E2GMer2hV5pJN7q4crrTss7kt4EecNt3Yf2LtGmn3oKdcvDj60U+UNwvudOzRdB0
RhNhorfdZA9DdaXm6lJhAQfUNZPCd7pSStudYHL0cyfN45OB+SoZqAOB9qTvGBN0
guOcD8hkRieKknppDNvanCGbOz/BqDRBt/GhwUHqQkDpCPYJafkNTbxGMGnrkN57
Tslfsu/ACaT3hC3Y4MZFINfakj1bH8H+F2jzEr/EYvveJ5GU896A4jTcbfRxcrhd
ioh0+N2hEfFQbPgX9zCpqqtX4nYphC+6ls/+yva3pGp+KgDHwbSHVhxv+CqhRVPO
QvvA46mOLmSioNRhAe7XBI5oOZkkCRuBcYuiqErB0z3c9ncn3tvFVJfycWIhpNRw
WiSS9Xc6LpMBuq2HZsG1G0seCe1fyLAaL/2pTSsX1LUCJRhJ2+IRChEfvx7EfU68
4L5d0EZz79lsFNNUInHlzwnunIE2BhK0Ux68htjYWESN9dFf17QfhxvCZ6Ho8Yd/
npggMviwnLiJoJ73/SdPfA3/63tGAh1rW1nZngpQjLPcgcqvht66v6us6jZzdM0i
TDSRztIriSRBEuokVM4yVb7V+ciu2be/zWCNAbUUMaFIj+JZgA2sECAOOnCUvCjK
5opAVyJvzkB1WJ4D6DsDLQVgT2Htzl02+Rci7SZutTTGlJnFPvfrjtW3o3TIXLEL
E86o0G41MqP3YjPzKK4nC826FsFMrNlWM5q6QGPFlyJzIxSNZqfxYZh3SWKIkW+M
40TihYVDgDjFssFOHbeqICW7zfnpkNc2IUxQdU0XCLJpBmp3F8ezQx5zCcdekk+m
DXAY1YRI3jwwZGPGxPXJFphUeg/dUJW52I9/7/W5ihdIsmSQEDrIUR5iMmC1zcTP
/HYXXo0crEu9WWMuD3OPV+FDXdQrB+gXUiYe3zYu29awkSBXQz5eZpYjQ1dJK6tC
18Fc5d9LEX02eeetNwA2IRvFhinfnSGOdkCXV4ldBA/AY7n76HLQKUTOO9ffCuAQ
BNw1XcgWpWuBv3nm063jYb3k12gCxB05iNRHFc37vVxn0NAAoZAM6vaJY2QuvyTG
sJ5UktmoXTZAl+1YF1pUK9hqZ4EL52u/1WwL5PQwswjjzEHzqy0Q2/DYifw0EoSf
2b500alhqNUCxXsFziOHxcT/YDPqPj6/QUtL+7s++jqj8/Yp1Wh4yYAk4eaZg4UB
MuVNzXUW/zq8kcYYbh7IYm8oRhS3YoPc0b9V8V7xiDEhycM5J5VvpkQmGsH5nbJl
7ryq82j4qZSBsIa3l9B9LvUs1U0Twtp8UFSs2OAoGfM9Oe7dBZyRLn5j5rx1b3sG
CUrC/Nyyy50cmKnPp8ye1GSvHrtqVajxboznPgLafKULumy9KG8UbxJR1B37DbWo
IMLw8yVagu3cusCLj/wZA+eAA92VQzqw8zMYkEmBxVSsRzjF3mHcPoT6H0h7dFv5
tWliLvjrmxVMATGX8UunV+VlKVeLSJpcC4vmdsRWhmi0q5TVSn1/styyKXV2dUMW
Mf3kWBp+dfE/MeYNyPX0+z7+ronexBL18cJNA6hcFRIK/yHq7pR1xFDgfGqa4BC4
J/j1X/xgh07qYeeKe7a9ss30gd2oKNfeGncj2w/qCDnBlJUcTjyDCZBbHqebjE1T
ve1CCoonX0cRL5rvEWDb5y3hLfSWplFnOupf15TgCVhcyI87F5YPp/cw2K+zslxO
+0EzixqD1fObKVUcBhrfhZJk1e8a1mePst0ovikLIeQuqxNFZ0cTKxuXIfZKZw/3
8JfvUHS9U5HxkwzNr4XQoCAGYymdnzjJMNGtDchbYqJalB9IKSGPitDqnpgfwRf4
V9f34W1BBu9KVSfdtgFP3pU4MdmiqKYnkYd3/Rgo458iu7f1N8Fzj//ZffAxukc1
iQOnR7MtYw9NuGVDX07bCymkEO5lo0Yh4R6j/djfbSnpJ+8oUW5dRp2XSaTelAu1
2tib3TwLTUyLrd6h0MWVBsoU0v7ueMQyY1/ZnvoUSH7VMrWczbAa+zs7QFIBwOnt
tulpxkQe5KczlUTLRZ7/Wb+VxaN12NhW7muyHbhS4o4/7J9iDdoMypsbcdTAqfKV
GejmVqI19PhHHJ/Pu8N38d3q2O1X6gy2C9t5QEjIoHj8v4Z1gJd4U6NarnX5BsMv
Xqmrw3r3olyr1Y/BsmzUQd2CWvGSS1Z4IrCXflhjR7EzhsaKO9oqjQ+do7LhFgCf
YNz61STlabtOpMcv0sKZfm1+ARDkYnJR6TvSFlHWRjf5dn+Q+cR/8cdZHulrznIR
8UmYUKox1EtOmqlWTbgLy1PwQ6LMOBiaiRjM9ynouNcpBimTndjjICQsqGl2t8T8
+vNbQkSPoaxcyziUOexlguFn46SqetEANh7DZaxE7rPqt14fWrgUscj/Y0xHt9pM
XH5toYLuEUhW0I7rq1UQLfOAHpo/AxNo8GMtpe7dy9CaKAKnxK4VknevpKSb95YM
SdLA92m0LoT8fSMio42SMNClRrnpqJxvQnrvsFVhRFu5AZHn2QYoI37I/bIlxXNl
Pj2ZWPRVBHzwzxbddMRupz6ijRTtPNIgwk0FaLiAyCq2O/3San/WiGZHWqZ5ZsW3
l9v5M1ZllBM+vaogWVrKJi14YrCDtysRLv+C5V2jMOf6XFNpPjlw8jq/306Mjggn
ntsBZfqdtIQ8L8YUoOKCvzmuprxCZPIZf6kaM0pe3RZcWIeH5LRHCnpbHxb7pinn
Dfc0qH6pnrlodkLmGgYLN8JR7PvPuHSdKeWg6xX2ULvoav+ty8C+Q+XTdLT4Qu2w
5HfZzFp5yuOAolVRFECbgIKjec1xB5Qbg1j+6FlwuIxrzJMHoCfgpWpk7yhUe8+j
BgFvFI/mYQ0NHbdeMkxcXym/h5AK9D/hRpSQbQULEQfv8iG07BbpY9fIp7cfUf7m
l9Wk9F2wMTEd64CEBaePAQmM+vOZVkTOwqzCFnrAVrFMdBPtG8lFTnWQwmxxwbxS
Hl6t7iazWt1SBCU5uJ8eTwKXVc6wnF4K+iD1p9BtX04CVEjaPeQCrm+nqiqReNPs
7ADHBmCodcY2WEm8WUrUNMTsepSqZr+K7A+BfqHjPd/NclbW76Uah+fRdYiTICap
P9CjTd0l/eRA8772vu8ePJE5LS/SUJGQ51i1tnB5Gp/HdXPhsfJ/vD2joi17vGu/
im5OTNM/cHV4bHkIdyLRr3p0ANPtRtxcR9qmF0XQETBcrI+Yr1VCwL6zRfrk+FKR
ji90sPnu/9/vcFXrtnxfBDeYcJNGFuc6uqpBCBBBCS0lhWCwqAumzFfHlwF8fHQx
enrEdlR3UaFtQnHtfjd3GcfB5Z0JHU0jbi15YnxIhd4SXSIfIwJ4FnGomJ0bcuf2
2AUgPTbY/IjSKAcL8Jr8/NghQIKrKzeyr+ir5pcTngf6S3gcY2IELBk1ka+L2vG1
k6ruxgj786Q02d1Amg6mT8yWO5Rju6Y+Vyph3UWIkDubEOEpcteTxOThzUY1bxrC
X9JvSQBnvKo9KhLuMIKqcmeCssDd/f9GjGqzXPksb/PFRPqABw4T6AhEgUg8kKep
8KkNsn59t/NmokhE/D01zRcEGx2a2aCiNmcDpXlvHA8V3vJOQG19JkX+aL1aMh81
h6Ilf5Lshz0n76OAUVVXJHPqF+St1G6NbXGlWtUA6VTd6MkMbopds3x3UE1nsqoK
3BALwk5uqXaKXYkmJutMqwB77JgqwwTzecybghdaOI+w57xm/H25Nukhz8r3thZi
ghspMicCeUChi6KSHQo7BHwPBgHWMuY6ZUsMdxTzv0FKgM5DWu/rtDDoffj2c14X
jItpJPs31IbX206L2rTnHmxn013PeJPkveacef2KbO6aB0BdIlb84gnmXg0u6CpR
z7fYKLOHrHSbeqehd7uYBE22kJur65d7IWQztRB+4MB2ritdl/3B4AD45b/LwvAW
6KNjGqmSWJQKygh3kR9GbC8XnrKpQFTFxIU9p1vyGk6tMBjRMNF+u+D3rBdtIrLl
vaWDQqJuJ0G+MeSCuuBMsZSTOwpFj2Ebonwsh91p934Y0xTsqthwHoc1fonkQQbi
fuRTChHbO4Fb4tinj5xZ2e5VovzomKf42U1oddcni+dqBzyyp76P6mTjTi2Efbgd
nIQToHbu3e8wkKbH1/tr4cHWXYJf3UV4ydvHGy//SPtDgOjiO6AiAex+IwGZmv8p
M+EZFiPaVOKUjaY/L+UiKWWM1oA+zK06y6Rz3qarhZdtApZ8zyS6/5C1daGmHb4q
KYfDqekJY3VPVn2InM8MBnQVAv09q5EfVua9mGAygh591twE8emndLdkhrRNt3t2
/iJUccG1ZNIP6eeo7H+UUep8V9M4ArSTnFv0Y06Xc5KbTLFpFCb+SAlozhwjEbcs
lA7UPjTMjoS8d/VFdfjgEy2L5DtM3vvuztn4LqSYqg4AJOkQckkpv6oc+WfFfYIs
j+crdofA/pt5ZxSyrhuY8orKFwG0rt7ZYNjaMpQ4BrGey1mTw9m2t4+9kuTgSioK
s2ZAzezq1M81YioYuQtK4FrjfqZloJhzL7A07OjEkmexwNiDOofhRtDTe5EAOhHt
T3LCbLL3mvTqw/yPCYy9Q9gkOby4j9uC88YgQb0+CaHQ4+TpFG5qxFLurYuQiFL6
pue2HngPgGxnUziXQUFRGjqbQfByQCLzen5h0mjTNL94rG/xshM/YaG5WLPSCGGu
Dlpn0jXPh38ozGI6NMMFRfV6wiBnY0KqIiFPylpejGdbbdFdPn4boZtHsFjg4l2h
PkrYW6neqQI6XO0INaVHZh06nf45XtKA4oa/JMJUTDcgyigSwCFc0WZevIH5xEna
Tp0jqYLG37uyQpFmAj29Se6Lll5SqEWWMasjI8UNx0P1yqe/fmrXQYUUv/6VHkbM
tVyFbgFQ/CBOpcAwG1y7jfdeji0PipGNTGbM3++sv6hV6Ls+728NXzUZ9iMiAwXq
aH7agJkgP9owTEaPLoPSXnk4wkHc8C71UlcscBuO3zAMxCYXkGAVhAFjT/ry1H9K
hUKQckKm/o7HqLEZ2pf6e6wlfbMHAA7OoDJ1wZvgwsHA3JGOcYni0EQ8JeHp7JwK
VXC9elWg2/+dy2099pM51UBT02JzB2q0ffz68jBflxZLb2lbuecNHqv/fH3hY2Ya
VinStsGfdoJppEclxzsI9epsljmsamebnSW+Hll0GZz6b/ivwEBM6ODtVH43ACF6
bAHUJTfUZRnqb0MZonG0GvEv1xC2UgYtgdHKdDOV0cRTL3Q2iyzdIeMFfPskl6ax
vBXx343CRo92/7+TzcfJfGzuLkSBlCQvc+cL2Ciz1shh7zjGaAe1oCgenBXeDMkY
XIcHevt2y9UooQJBWdt5oyCu+2My6v16Euz6/Mlk46PQhlWXooeiB4UOMy9qMi5F
dhkKlBZE5LENwHwWJLk/czN/wrPzYkUN4c57gST8OSikTDvblJoT+5//Li4WRROE
sOf+YVFpZSwRaEWWohDeSbUazhQGdRHOthwWhvrf+H5Pq07QPfcHGt7QBUL3nTe0
sBmIi28tcYzYiBCPkmdBkwb+MAPwyjiyPWw8b1AZN8wQ0cjyug7dYmsT+yjeClhF
BfUsRQuKXGc0NX2yLq0p60FM4KwpeA9au67f66aa4Ab6oMz8AlR35jrkKYK6lwkE
MYnuMk0PcoHRArasXUl6RrGEq8lXcSb+7K84rowKe5ai/pQTHZ+mcAgT+UPHecsG
kSRPfV7e5U30Ikvir8VZCRue4UQT8SfihTnKFeU2w4Vs99xjr3ffl3P2wQ9nvnFk
h+N2z8TBPmRXUWGvj1NtP7qZ4mslnanqp41WCJl5T5fKkhmkKRWK3rHX52FFlREr
5GSUOartoaXQOKFd8Rx/B2JT6VgUM2loCPRm68v4SNh5NY5Fwurg7qIGFgw3tV6x
vOfICa6Uui2t+SJH/HP69Z+MTSugnA3pufMvuNLSjOW1lXaG9kllGHEe7xWKMc4Q
ihBlkipplhxww6RyFZ0iNXzVa13Kui8WFCiGOhr9u5LG3Lpybs5xT01p8e2wnuX3
L7UVeXl5uiihTj8C65PtJGFDBLXhLkKlTFxwy8ZzBw9HMDqS0X5r0AlScD65LTzc
qSdOushYb2FsUJqNlF76hgKvykwdTXJzoFrYOmoK9TmFJRU4UaNWEEGGEbTDvsm3
+eC/7ya5CGAoeZKEmKV5avLo/TFSAmTVwsrLpaQCaO04RsRIz3wI/FwhMMMa7j1i
UfGmaSGRG2ePZrCEToHBPAahyaF09m6M5SBoFuWIz089k83fCVHbMqFfpYoF93BB
DAMN1wXPXEScMZZE7nHcoZ1eJQwqJ/cTxWtNreO9d5al7JOAZEKl7ba6BQ3/MqIa
bApnBBQ5WzVp6dvoJGnF2vHPUz3HxkAWdcxTdzVsy/8b+aSDS4R09+shqOYVq3pt
fawuLSCpklLLTrXHyLoZQUOKfSGIyr2gAp3ITAMK7Rqg14MmVW/InIqgiooGu6Dv
TrWRNJ1l7/tci+IFnrEtiM84/zzpoO5GjzYnmiO3A/XacyhH/wHhR/2tTqTTSr3O
mWf5pr8D9E48MYz+J1u72NuyTE6YYMQk7u38rnidOXObTEKL7wGxoQjCk1f6JIOe
ki0UTOpouOtSk9YESoGsG7V1GY2YrcypW/THLU8tgy1mvwMB9DFk91OC36m4lIUU
ABZfNxHsd2g6LC0qlRHJqm5g7v/qfHnI6icFgN0CT7777axpaVBGNB0UFWFfuQPI
LlKDn4G2EUyvnIOvOp+79flpDcsLo3pXbEOW8WWg/+Ugx0xXQQ3HoSPTYrwZsEHD
0DU3X0cBVjDe5VNQ/U8AdEHkkYFBKX01eX9PGs5DpHKELvFRvXBgpCRlTdpo0P1E
N+avhhfbEgz/RRZKeDig+KRc7M2zqQTRDE0E1kH98KMsCtUxEYEVNWu5oRI3pvjr
piYy/tpEGEpT+DWISh5h/2rdgWcECgk9uhY1WeNKWAUIrOLj4iBE18GKuxJcMYLu
yZiRNTgECfuUC++KfPOetD8qjmoPDDp9E21OHUF8zXnDTihqDRaxW7hjrJ5xA4Hf
h+hyryxNBBHQdW0RPdIDi3AuGJcdPnUJRwPYvbhfpqo1jMDBWGgbY+vUNdfG/ze1
18YtBRP92phfpHzdawabq9medErWvdKCP7AtWIKiOfRkXfzsz0R/U1mUjdnkiGM8
4r7payz9OIsdpHXmPDMLFZqA+VIsK/QW3fZGWYTfKqzTRTPyHUKzNhyaFCZGNK/4
K8x22sfvdkz2gQehMAbuEN5CYYRG1wMbT7lbeQ4zDAg0gYWgQfSnv/fM+whuRwoT
ClFKHrGFCYoanmUpVH7zCzG44e9sHzGU9vKagj7I4Otz2Zw33lQi3KObVijnrYFV
dzOv3L2V8+3Xa+jomyTkJAfnb6gu/+G9helaI4qsL1l111oa3wF20NjNpy9SVnGa
UbVPdc9BlJW7Drp/qfKldJ50o5usL4IZIeSUZyAGvyv9gWjJJYqZAQq5sm5eDVrO
kfM1Rqge+BDHYzSS++o3DC/Kupx9GBPtfg2jp0qq1HJwmms39NhS8+ff2rkQrTJB
e34gkQ210hmNg9voc9jIztzCfXxqBxe4eFMORGbisNaDCDqMAUJE07DmJrvlyuXL
OW0A9Zb5XRroTrGJP2dZ6a72LdPdRQLNVWej5Fdt4GdC2Ao+cmm2hvANJSduuZJf
DupDnEEr6qjAWLii2QL+PbkWD4v4tJ/co5JhtKHPsk3nA2Hghz8Djng5mwgGrwGa
tG4w4zVbleVO6qypf4cd1MJxBEhfftSYO23nWOPQke8TwXRS61w+rB0hpVrOMJLK
dBCw6M6YhdTSsOmn3LRGMjDdHVoD++UvTB8CX+4q2x1Vab6XnNLxA4o8L0dT+WRL
j4tbctRXGy/XwemFuyHZauhxB5gCQAEs2oDtRvDbRU+PCbsxDEfdftHby4L+10M3
k2LGgHyB9k2zA9Gb5wbret3b/+SiIIQmxRoifTwytf459icB80FSckH7N9cgU8qj
IOuqnPWV+LSaYJ0KxLoOG3evXs5MYG2LrYFzquPq0VYgUZP8jiaZXWyVdCWbryeo
TleYNvD1LouoALO6Fl5uzzftVLgb3mRC5yaRYQwB8i4g0Dkfoz/fQPTvAlENFFF4
D+jbbsoMPYpgd3ZIx5G1EcPqWLkcgwI+oP5V1hPVDrUwcITaduiFjIu3TShWHnrK
xAa70qF8ksYDcGfJFzC4k8Pq1rwY6oHI34Z8KkcMdTIzK4KGW/ag/pV+wYGUC2Ve
qoVniSZk7HWSSW/qUMY8kPBvWHCI7K6S2gExesksGm1MTRDhZ/L5k+4lQ8DooHxP
jtb1MqGiYnhEA9BOdWneT4e+Bz1NEYTwlxSCrkNu7/152/9cw/vwQRXjZyg0wUd1
F/pYQvUbeHefKzzpN7h93jqSuf0p2qq2bA5eSCTK4iltpAz/cIaVFFzzn2xCALiU
bIUn6OjmZ6xHbMIjAQ7eeZp7QmcmrqB1au+UxmnVE/kWQ4pFo1DC5NbwVrSCXwbs
+iY049f8Ab6NG3rfBHFDWXEi1zZrvIC43GvGqiOy/O0QXOEtaXPll+YHx9V4N4iS
WFMpz5Kk9DT39OeyY3dxdl5d3MwpBLevSTWLykUtCEc8RVJahQG94n/A6XIiQnKq
AVesmczsz7dbQcv5Y7Vv9kv+A3HZ13bTgIfOeaUMAbESJUXru+q6cl0nlTVmfVZJ
nKb8zY57gYKU+1ra1BCerYah8nO24p2KuOI3Ih5C6T6hSjzhkTKmwqqGAV9KCaFv
5IXCtJISSHG2Bc9tNkkePopYuBWZeWHbk6HQ7QKZkVt1gOybFdnYtv5mclNDSn4p
5jX8Ty86u2q1s7yVAGHKbbKCkoHK9jZilkfRnCBH/mdZNzCtqlc6ai2lUJ4vWOJD
n7qjraZO4RbbWCfxDTbXWaH0YIislWflghCKlwoYyoz766euYJECnwsz4T0o0ZSd
bgPs13qQdjX2OITSJWv6jKytxVdiudwtnr2J6sZPLsfk++97rgITzzh3Ac+TFG0B
FJYX4/fDei/SsAr0FXEZRyOyOeGjJjNU/1hop3KfZoUQiHgIr3gbTV49kBzkbG2L
CKhZdlgUQA8FHSu+t09L0x4IS5YqPp2Gx/q7AqnP7Kdm6tKYaByhNQA/Wm/1oUD5
te7TPG6XmVHmqke1FLIBBos5XK4pbHV7geAYqI80qpkIAEbeZuxkqaCmlKiyVyYH
p5QhKt4VqbRRViNqIExc3h+XhNm2ZXn9BFbXA32jpKsTQ5LADbRXFi6xvf6gejCN
RPqiCs09VkbDYIXNz+w2yQ7x/ZYybFDneb2h0Nn2wjabSaE7J4MjODjp397UhlcM
GnzkLdDaoDGx6pDpAdyv4aUNcLnDm1yqoUqdpoV5gTxG7hkamHIeYqtP5DHCINBT
4sR6gV4o6QIQEWnXLdcE9hhrfA4lERwnbtU5E9zXzbPDoU18waQocPR3RutKeEFp
VILOVe8psVfcm/pfD2ocoETNdgWJ3RaxqkA01M6N/tWiZEySvxVzDd4c/syAnNXQ
mixWcJaaIHUHu9K6aTZCr+SjpBro1RyrN/EDfPsaGqR6RROfDHOdXG2d5/y7y1qD
cP8/peC2H+4tMRUCB+mYQoB15rEbbNfAgCRCd08i2BH2gS8o6N5MoP4QvgL56eSC
o4XcJ0mMd6gO9zlua11zf01wVNYL5yb2tRxPGeurWM5Ud6O8GgzSUbPqsG5y+KyD
hkC1rKm/LTn51CgfGgEizjJPFyU/3WYKgBWFn7v99i/K+YaEaNTl6Qc6Jqhe+R+0
7bfsUTuyp5yo/D7szJo6alyOQTwX6c4z4UlX9kWdjLNJbtJVYHLJSS93/1FaheJC
y/6KSzCNXMBsj6qWFSxtM/KedCgkCwaY5BQRXGzd8+HrdnZZ2kclwLv0CEOzy1LN
DmT7hFCeSRdDwTUi67OvOAB8fn/jQnadTworzxEtkRoK8SeJwgk+vihewH/1VeWY
tphiTr4386+a4Yv1NYiQJFw2C9u+NFZVB45mk3vFfHFTrT2a3lu0+BjXTBueZWc5
8n4XoqvLy4G2VlGx5iEYh91asg5J3SWFqa8tbcmsMUWbTI/hNAc/7SQob2UiI8ip
MVMtw3dckvuTr+3CZfVpocluVq50Aix4WraYV5GdgWJ/koIpgCV1NV+ZyL6m7bkx
ZS+qXOtdsynX6EoK5pBAx20mxvINaEOPWZRLYXCMEFcpaAcI5qgVKVI7gCoiEKic
1GDsPx9c6YrtaXCANwYCqrQa6YPzF6JQKzHLwUUBnmoIJYflWorNufrHcnxKQZUX
eZMeE9aDNAFKrZCuo+Z+gBENKYlYAxIhPGwB80ReP3yU/Il2/1F4Z06vlz7ikFJq
HIwOz5ERcSEhzOeJNcJgs1qj2kfg/odrbTgXyIEvR9f74XjkW8sMHLKUYHlWn/hV
5ggP4UxGXM2ZIPhfs3c/obh5r7ee+yZBr1Gv6e9+1zGn939+x8+Su3ModmigWL3/
89ZSTJtyzuICcQ4WFvCdt8LZyP8edSUz3i4g5sSAfrZYJQiD00XpYpJ+rB5Pla9m
ptnVjdZe3rqFmxLtbNjNh0qpc2sig6kDKaF2hJ4FSZWhaYda7KenyX71jHUXuS29
fnO78TxCvjT0AT+tJRaqjm3BJEfnErlnyi8XnsQji2jMrBH85KalITNUJLoaHTh4
4wqqCYgHlJPvVqhwFTG652p8ZfV5ByXizmWyLlVoIO99sFizF+9K5xY2uB5XyqbU
/q6LdXRLVh8Yb9f1BCzVTFYx67nTO+ad2Qi+gjIngthULbSNpTZNsw4LkhzLRRQr
Y3v0+vKMjwpIq3Sppb9sYG1dOkz4B0UOeWmEGUOnAp2MTMO/wdtOOVZGEq/pzcJ9
+gHGsm69CR8iEzB/PLWmWpEWW1kLBoZxZygQcaw3Fwkso11B2lZwgPZqHNTz4W8T
GWpppDZ8A7AWqQiWgn6yXh/Zl7334E+bRN5+PwedoS+VRJlMSkpq+wn+nUx6m/oe
luRnuFH/+Ti49Q05Cb1t7z+r2BsOM8Yqpa9A2gcge+g0Bz/c1y7gDS5ChZSmz7Hc
FqZ7DPe2RXqCYlQUhddNSLHEXTahJBx97wZfx5goDwdlW7T89tiO552IWUK1E8ri
LlLpjdS2EdQ/izvqYobgB9//rw/3aDRH1Gx3xIdP3+cZ4r3pklkfpFu/KgL1LUNP
9c4Rzxbio23mPldbTfhUVd7Hoq15kdvvZKv3OlfvbQ9ek0vTour3qw4EsGqM8QNX
QWaHl5dYAI931oAuLJjkEklfUhgWB6Rh1m/oobby8EJ86ucywqaixLk2vP54qgpT
ZYMvOKcMtQ2KfBcMkU9MkD7ok8N4czS7ImXNiW09AgMvJzgU1fpgW9mTLgqefrnJ
xjd/IC3ep+limgi3FcyvH+GMf02Bax51xvl+5Kv8VUhRBnhH8wVQHTcxKFXuWV8g
60ZJHIBmzjf91GWKlWywnFMBBadTBSBn9AKMwsvmvpso+SDFddI2jdFwMRqEyUXi
haafyF/3E2WPpKF3T3HhTTLjtmwCJZ2bvXIq6koWFRGo9G7wOXwwih1jzfHKZeYG
86DExMAKNN4PPv/qxnmj+SiDij/hNFbany+C1SFjF9RqUuzmYlgo2iVrs+Vgr3MK
c3EQK0U1uzmnq0RcriwyEcC0AIYfhzqu7OhEbm0ct191Ya4ZJqwQfMKx+FqLeEVy
M9nS4NV7raj6RqvNLnReXh8xhWVpYA+UVSAL2fYrHFdlmbn9hY94WkAf4yhkEKiR
jGMGyoU5N/2KqZR60WsztYuw1WGXRTla761judVqvV27CaRfs4zXTeJ0wcT194E+
u0Nqf8OETKDdW60H60mN110pSuso5ZwVpufdXMuL7N59ve1aC+gfAdP5QhYDJP3W
sm6Hs2HwvAYXfraLt+5vay3P3ySE83AgJr6zudFTEgROzoaojcx05kXP0XYdzc6C
YzXycgasakJp+8eytSex5doGxzzEbiTMhqNGy6FmAFzUhqORCGQyRzp51+H4trNo
TSsSAHJKHDR1zbOI9Ex/D3sIVAJ/A/5Ga8dmz6xrisFql4/nVCRIGXRRyzTJvZfk
SIlbbkxue6+/XY4+2JIGxf9+WlVRIe+zzEkGvL65ox/N39XwnsTsfSmaHHZQDFNm
IP6L0raVksfIkBWqoC4qh/b9oV8U9cz6a0BISSmMggHNRaEqJpkT9hha+dHs2lsf
jLSTqeqa1GXL9vAC8CuWlIu6Ud9n0OaVg13jROz1SMNV4bpxkHRrCdcG3ymHAOln
cKqqagR7rUxlcM5tHmj1HGF2TxZt/R3z6Nad8z4r6Z3RaeGxhEnF2GVhs0f/nPPB
3f6OfC9bLZTsp8TFHW64/fJnm7H2wkYfj0XEeqFcGr8dxFxKFBkaWeqLxYF/7zel
30pnXey7bxMmsZCX7lRmiMhHjmbxOgruj9BgPgBMDuzWk8wNlUO/Vj8yMWErA/jr
lVz+LMWVVZZ3gowJB/fz3rsKrG4PGNZHHcnOXRtgOroI7w0wTmQBLtkvJFun9sHU
tZ0cRNXTqz/+lyz9XXeAlopTphbpPd5Eb6icvYyaAMd43HxJzSbx2I9c/LWK/kDF
ytqxq7JOwRSGnd5MaRjo/jEL63K8Dtaczma0jkFf5MUtwXpehf29znbDD0rSuJJv
ZgJ4pwkXq9Akmykb2p6KH8pLQMdGmv8Uzx27xlGMf9GysILZRiIggZGTYa+0auov
jRmoSG4/ebwC+5DsOzXZ13T+kVjuowC7HQvIMbciVDgkYvTdzdRMcEzryJ5md3cB
aSE31BiBDbt9SgncRo2roKnm60DflbQCjxLzziR0srp561FJk34hdfij0/cxEgKt
9Wr+7qh4O5nWjSAOgD855V9aWONInNalb8EhE5vvejYLvxQq9iyKkMiySOBwh76R
0pDjdGp3adP4GA/P6ydSLypW1nbhVjw3ojMQje0NoB8Dj+d/OtLYlNnn66GTXn/5
J6yo2Xg7Nn4ql2HdgvxuwLWhjkHi8JS2VIfDqFxbb7ROpcGO5ExQOp3kynPmbwWX
Wto1fw1geAtMwQ7CJkQEJHwrFv93nqCBAEIUVeOT3JDdd+IvQeaUJZ0VT0nexZx+
RIaeC7fFNszNYWjmhQcQeTVifbr9D6nyy7T7ll2lnSR+jzpGab32X9kwSINzpoSi
tqcsEBWYZtcIFgRLXmpAWgfXIlti0AlmXbOeqYzFNqiRFoqeZr+lFbLg6UUrDmQx
z5nm8bxSQRxn29L/Up0A6so09B6T64buVg17PYu0C/IJ2TnVx/96nE1YcmsMZaDz
c+YXwJD+HVLUaP5En91NGtx5oJ+GvEOSmgZMtyNb27tjVrBWS0VtJmOtO/yvZJAM
Is9B1jD2qS0WNoEGWvi/ft+eWPZaFkfUXjy3l3eTblTQAncHnXz+1gT6mC8DaA+e
ZN8jQBkwUmS6nJxqWDR+2DNSPLE5DQbuEWec/vv3vjeTKsLttXINcQY4sK2z+ni8
DAWMj6SQ8utkx3sxLNkyD4u2Ugwr5k7EmmLqO641dramm92erP5uPpnh4Pc/0zXZ
9s9mPxEduyTQzhAA5htJWwkA9EFTTwiipOwfULo9FPAJCsS8yCjyFLAgxxlykzJ0
jSuw8hdVlZHIQe+lU23xoG+xqZA3yXpsVO4PtkNsgCxIz+SMCKb7E0lZ1R7Mps3G
aM9GLBTVrfhhWtIVjwS7NNxVW8TIjMMNP7jM+WgbWVzhs8P3AJ9hUuzE/XoGMbsT
HibOVSPNUuo1QJrPNWOeCLA9w1AxiugodB/IaRQDXBDcM/8kZPkSaYnNj7QXVh50
+V46gRQJlz7FzxIqowKpa17/oMYjtPRCHRfM7ax+gzY30nFtT5Or15zPcmBZyyw9
+9xOkJcC1u9F358L2hmqkpV1fiQINtCv7n9Ijh+zEdxT7BgV36o731IqsHrdybed
wlw386T3rt1F9kfqAP0VqgYw78wZf/xl885OjquteqqK2gJOXYkhbtMg0F5UEaRR
0vdzhey4jzzYBQm+Kz678esPJ6MkBDmQuwTE+Oz9cKEyCfQiXfYGeh1g0HQ2Xbbg
0I4jTOi3o2JgM4VxUm5nGEScZc2/hkII0ttrjZbHYmvbG1PnlcrEemJJSAHyOwn8
OdsIDIzLMcNpwCnsEJEgIXqqDwvg7Eho1yE8PkvTkKlgEPDb+y7lw62T2KHZfaot
zWRnR4Yw7KuS2Vlifwze4Tf/2amddsx+LEPpQwsxtYaH4EPmJ3KzDRX0MDWVJfMj
CIHPzuTaK0n52m6QP+vdoPxiw1Oo5US66mbBDq0FNtRwsvaYGXmGmmKagUmNTMs+
b5xiZMzHHUJsnqsWXhIINgf68wddhk1kUCkapFLSde13VJOabXiUigPZxt7ivx04
b9hqYte7UIL8vzZkrqkaQWAopwKWlKIANUYS4TF+1SK+GDvIrkcH0ZgwfRkma3Yl
HovV7H9AN6l5dDE+POpK/YGrkyOyylGSAgtKb4zuJ2zRy6xE19rBnvLz/ztnv6x+
IqntzA2E5NH9jKTKPM7XJ6Skghtwv93xgPnCxcZunHPBxaBIK22Xy068DJoYbYSu
skOPHv5am/Ty5GqZGPHkFibeJUIdpLbuknCyGAhMuzm+knVhqGKiW8GzpbUwkQY4
J0BYlUqLZ6IKHUqKx3CaGYB4urz7sf6c1rnb9p+65bUS/+ZbRgS7Eql9QCy9uHip
BiyF+Iaz+2kMweSdiPzQmPvTjljU1n/siDRnyMNChVco5i1VmZ7qCL2ZUi/uDO5a
r9eJXMnyRUKR5XjjcV6ZAcXEMoYf68q+8au7LjAMa6wv+6pFl6WFV2F0KGYL6yZR
Bdp9j7f61mZwww4gIE7q6CQitjvzplY548KQzXhDbG7X11ZS1ticxbj+K8J1w3Di
bJYXe4DLLQwA8oNK7Vi1EAFaSRSMnL9q5otalrWX7YGWsdO9Ps52ZsIOrgGPPre2
FcUGNIUBK4J9F0YM/X0QNmyvgotWO+SZG3Jpviw5FTWcdhh/5wRWs5h/hMzrOYDP
77PmhfLFsRrvXEsFhC3cwHkIlVAumyYSr0M7Yu8l6F7+mN1CWwHTbzBzQ6RQg9WX
6Wj10yc+CbLrlqgP2LVTx3YLwWJ5+YA2oxZxA83OkNMrCDSZ4DzWO0yWZFEg0n/G
5yQst+g6SGRQgoFqXfPqWvXRd07Tahqpdf4j7gyA45aMy2qnVGbMSYTO9ZFwkxf3
Nfc3xcGZxR+uHhnzveaR/76hlutmQ8EGcpm4v7KpdI8M3IDQYTYBcLx4uxiNHK7L
q0TOxgVQAlsdHbvRHL0E372fVVPtOWBBHLBlax0jGsRd+imcglrH5QcgBuinPdsJ
V5P93gPY+CYC2WC0Z77m8/K0ewI0obEnDNOH5TUGIxAGBOJRdbhClO6LWphk3q9p
DSDIcxgVwNzNXg8ZEtoi03wbyllzPQbVpqB96oL0WHQo7l/YsSVIF694xa5LlgTj
HuX5MziAX+ULKP1v4BUSLvIvFyras7LcH3QTh191qia45qJPWyWGq4yqPWpxXVAW
T5KTFbD6fYYzD0RKclaTV9QeNR8GYO/L5KHpvIPviwy2+7EyHLveZCOhCDvOWJYP
+LSj+7qNOIRGdJAAiGgmFBHnQrJg9aBaDRpvENNNbW28DYJG1IcWwLNG9F/hJAjy
Sciw+WYEwloewRGUcT93znoleEwK6V1RIq3Y+EKSmfpduFKzkLivtgwVdYFjhX00
ZecrtoGpY85G/swpg5zf1cAsLzppAoVnGeUBQi+OJ/048eU291aIb1ucDLZcp364
/z5A6yEOWbzMjYuXi26M3RQdUJJ6XApa+TZx6pdZBiAsTWvlc/3UJG1j6CFrgNyE
QyKtZq2bZ0KViteW5+O6dGuwnoQqmAmUGuov9Nvbfn6z+xXmUDhFbwbmY0Gvexoj
HrvMMxo6qNYPkIEcpXTw3VLU1avYKG2oePfmuSqpfvBZHjOzV6S2dl18rgqarPZJ
+ma6sGmklG4soHj8nKAobQt4omkehpixyEBQCUeima2Z3znOOQJ0LTP3qCUucNgS
6QeJyA1POWrYD7y7LVwDcuv/KUHMCmftO/OMh+WqjhwWgct5pRySxSB2kl3SfSt5
+eMJy+M+gNJrgsq/SkDn66cEwa5RSEurvrA3grjUpN4FnXAaYGu+Z7FWO4FHyzV6
AqW35clN2hLU0kvoafyfUjyGIbzWirnh67Lc9vLW7DZZJxMhXz+AspT9OV/ar5GO
OXRjTNPd+7ELcqL4DdaFiWrRbNnFcJoL1N+vB+lbDCoo6tSlhadd5rovePzQ0Cjt
MefmUJaZ69dsdltIZwnxeDPHbYz4jSSTRRN9fEKGi1nnlbWOVwUSLcf8lnY1fzKO
eNg+Pd7nVE9spBQkkgPxi10Z3VYrxpqDuN4cwcA3Yc6JkzfoaHkZOClPpeOYd3x0
FlKqhPIWIto5SXnDDcvon1AI4rE1llRGY24TbV/apTlRRmupG9aUVF/yeQAfhzyg
yyN3aL2vGqK+nSa21s43MbDbr9uluoE+8z5ExbLzOwKmfRcsDF8pdRfgNhpjPV4S
P0KDdgRSSLib1CrwMQYyGT0yBze5NIHUn/B6fFhd+6coyF55EKhUfwy+KhR9/ZzD
0K4Iq6JD8dqL70dOBWyvYl38IhE7aXLLOUHIYGOCpUdLt+gwhveYqwwyVvb+z3Rc
0T7D5tcuwYFFJhSFzMHyHy1QgyuSli2tv+7Z/6q+oJnrjoV0Lrsr6zvrfEdc14Hy
X0twlr5M31L5pOQqrPsmzTtK6vEkfi3I/WLo8793C5nuFmqQ+Rit52N/RvPwNn5+
7WBwvIBHVgLMYUk2qxrHMFKD96kvgMy3dzuCNmsflxNfitNSJPUvaaGANtbp90rW
QTpoKVeRu+enkXELvmOzkmpRxRAZwE0qLeikRsU8mNlrmmTUXsH9mLvuepSI5rT3
9E1F96nzwvwSaRRYIGJTVz0JyiiSWZLiqIdwJ6DmDGKvCHsvhDCbV8pNAQj3QFpQ
SPiZ/dbkdMszWVSdkgO3UyyCJHlja7FXlIc1JOTBoAKpGuGTLDlqwv2t6s0kltKx
oogwbm5dYc5dexvKmykQA0jxkVrOq60LRI3cy9mwzLlFG415jw6cXih1CFCyUV3Y
tkv7Ws82ly7AV86gP1Btx+b81y1nK2Qjvv0dOKLggwGfxfynYBfdB32d/ScAwPSy
3H7WY+OClz4BHZqZmGor4vqU+dCeKvVJ4zqCIoXSFh0Iuk9nfVnnTe3uOdPeESCo
vw2p1BMUAF/ksYpNNl2g5nIA2hBpHi4hFcuegUl93wvG/A7GjhU+rgpZxIRE87fA
gtfRMzQ4euuQVO4peHPQJaEyHWI0ZdFBUc8Xa0C56qMu5Qtg+E4RA8vUSi2AuNRB
DqilRA5PVo5y3OMUuZuDoTqBc1dtvnb/QIRO6SQObCXAydaawAzHrKxRi82dMwkN
WuI87UwuGSzGTpq/qCZxtxB5IygLUKQJjPdbCGkmDO5Jvgb0bcQoqidZBFUsG/Hh
pTrzmP6PeCRaXER+aIJefYu02NG9tAb0MjCNW1SRqHqDbPmSLqMf22m0Hi3XKXta
WZm4p8L1akxVJBDOpC6YC/UZGKBg5k07SlJdLwvDZtmK2T9r+W2s6W+1oMTT33cC
wtRH3F/NKuv1s1FqD57PXxMt23zVLtSITJucB2a8OIKw+oZ0on2JrL3x5z5iqeRE
23oVR15tAXHZPTNYS6/+Z6pIQGMhnHvPFUrIXBC8eKxkm9WxxR+FSXJyksRLydCR
CQwiwKqkjhH4NYsTRhqDpvzsrcWpNGEIroTfKcvCOrjqInS2vykxs4WsNi3onQFD
S+RMIfoc6kjplQTLDX9LhAFkJExNcvHQEPKcbsUkPJ34F7RY48R013o4O5fYEMK+
BD0R1HQouLa/4fZ0NBYMHb+tmTehbk1oz11Bw7ZJbxPRS5Fhbm4IsqJbSarqFk+B
Lx4QT068DMV5nq8vLMN2BNhT1nmD7S/ZZTqmcre3zFMoewoIpaZzI1yGzFVVxC9J
wM6ETGBSOSyZPhk0nRROn2YuuxIcJpCBd3IgB4UqFPErVPZghlhXHELCw7x3/2kA
dWtymBH32bEwcHaJLVrOAIdd4tqJ9vO6e8Fvdjd5QUopzIvH4zmR4FCDJrzjg/Ws
kkljJcNojGcPZnkeXetTI1vl9hiTcMOYgplCnn1q0ck+11WH7TSz11zDT2U/vvMO
lO43rTUzYoT0d3R1lQ86+AkfT0g6NKpAqi8y2MSrf7pKYHszD3ld4lTR7gYd2/k8
/Vbe7Vl8Mfs55qYVGeObZcMKAWFwaOjce4FsEafRYLn48cf0q0E9MjSCKPMk66SP
rWQoS5fja8QTkSq+wmQqBCmJUeauri5PznRjLY54wI5ANoiHKJHrf5feVOCcmGK1
+zi3oMW1s8duXuApsD96cuxYwNtpUkHSjlagUp4epKG6xu0Eh2zHFYX2xgbaMR4m
lMXme5rEi4MEqSevGA1TMEvjd8eFGyjFN/vpni/hQVTu2Gc06gWA0v4bHbAsj/cE
LDkMt3LbJBupnllAnoX/Nea+Qfo8mUPBuYCIoAsSXRAHMxdAkG4wu994ELpjfvSk
ngQ/jVs5Bs3vSezNzP85FcRziLW0kmWVzn8KP84Nnx5tOtXiUf7qxZjZOryXdPsa
Si4HdBS5kXuRum+rQan2Jr7rUVocsa5BfZWjHxKQigjqtJSIXM+jEIECGH34Br3Z
gI1F8IfcQqtATz/5K2iXoJkO6L7pYpDl1ff+xaghaOvTrIEX8vUz3tQZe1BZIEUw
juMh80hgojXb0mHfEVSLRxtTBGd0zpS0Gqu5qpkXT/O7hvXP5vIbAmxqfWVhAfNr
Z6t2FUuYBeT7o+Hz2ZUFkpWCvPqI3KyDUmIfjL/IBAansRohYcmVKEiuD9C9p5tM
8gj5SHvSzN0DVc2ho3ETp3TFFuWB+O7RH+f1Q+eT0crgnN8CVqOE7YzfQqgxWd7K
3WFuhMlo59Bcj1u2gkuS9I4WEx4GnRBC4x6+Pgnvv1Fu8HKoLPJ0b4NcB7R+cW9c
7a5votxZY902vTCiG1wRjQZGNseJnlrgVuo3fyXPXUIRGiv5iGD2mp6x8fw2Z5rB
8RaqA4Ihi7/nls4HMfUmZ4zrm5FnLB6QGCsiCZ15DjO8rfmF021NPXAgftGhQWM6
vtE86he74eh3a4BwXfDj0mY9oLccIOqBlM4koIfnu2oYBV6Gk4GWyJWpHy+kkCJZ
LrbONtXe8GFaBr4p7ev+tF1VCQ4jPjn5FOe/mjFqe8u8Womw2GFE0Lq5ruJcfLGO
+rR8NTB/Spte4VFUYzG0Vi5YKkFTrzGPIn/kcg+d+Ymx3kZBp06SL4dtz5EwJd5Q
KRh7TzYHv5xB+AlPynD4KdsNCIQUfEw357x9H+I9nqw0pYaMXMpyGYzEttISsaF+
Dk3KptlCok0bLRzhHwCWoehaVB6YOG1jU4h1fDFrzSTDKguCVZrk2ruC7xwcCd6X
4umH8Lvxmhk2Ep/+Gwc2jxAo2Regw5xzcDUaS5HB1sm2Y24QZwroh5hDmUF9LNIK
o7sNDw1Tv8igU4m7yvXmvFWObGTj6TXo3SiSCPvb5LOO2ICgSyzDGeRlMeFqlFnb
aP3idMGNKIF4/FziM2vDaa/h+nzrK1bx2FMzGiXzCiJN8swNAf4bqu8GXLQP5DR1
RMfu+iYJS0RI3sPj52qz/jeG92hzzMLdrfVIET57n+feVcldqBO3e4ZaXbohBnKU
A6PlXiwj4ezYyuYpVL/oXUm4FoTldgAidZl0oOynYqLQySRBZOGEokLCWMQcsZtG
lvyTpinEhOPdVsfmruQmM287QD/yEGbKeJofCAQEG6n+Oau6oQLNPdCbSFb1pVj8
viFtF4eCBV4BxEm3RvxXyCPJ/RRpEVEZnqJPQL0/9tFIBjv452xSoOZLTaR0kK9w
UVUSchU8hpHdXwv3TR+bXRXOz4JkGMDtoGJ6rVC++jqLUfG/ScP/7RrZByi8WRzT
Hep3BHZ8DCg4BZP5X1mICgXFsGP3dPMDrcHPweiHK+7yI39LEfjmWoLbP17FAvy9
98jkk5xAv0gCUUAULkW9caYK3VBHwJyHuZ3Fr31hWI1m2MKYO9BIJfnZ3WhDVoTc
gjf/zRSsTbrTcQE7tdEoGV3HaCJ0B77Y8W/AxEXCQEC5r7XqhQL8b/Ky1ZwcJQJf
22o6XJLIUxskeohCcUcjyCQUIrYbBlEXYvDO61dk0XPgfrl6nMlJtoyMEHABlwqJ
8aAM7MGEvbqXilt94izVcF3EXpzp0lqlbzaDktJr5L6wmx/COoJJlWLyc1bZQBlF
y41GJtMGAELKL+KdvhA9huzYw3IXrcZ9M0Sm9iN+ql9OU45LKp3jT8u9XBQ4FGWK
UN/fAi8Dzkr8jF7rAsQXo69bQJUzMJvcXpSVhtc+JQFVTQrQ/2flOVcPDuqW7waQ
L233j/vzvj8tj+T9WYrr/yXtyv7urqbj6EZkUg3tET1MU2xdYz4JwEVediBnQRhz
qIWRcNniDjVHziDOyXD6WN7QjoctMZ1r8uEGKvPbGvJ08qyXYwjc72Kh2aVxLOxy
OW3hZ8CbTv6xq2//Qj56OndaExDL36zrD+Yy+CT9hZBpb3+SmoHlR3qREBVTmCjL
ZAx95T99n9I27k1tCBsc5koa0kzfwstPAMKqn/SUkwlHNFqJa3hL8ArB+72DTxRx
ljR9zBi20sjRB1k5An4ttCRgHNaN8DlzbfIFKyqDkwh+XWJ/jm8ENSi8lyFhQCrt
/irBdfTm5lcki7TIJQc/xYw5j2k++FR7E0ahL9RV5rgHIvwKx2pB/D62fTn0CK0v
CEu+oWRZEIaE+/FgwQlTY/hG+vf2xOWLr9/4bCWyp1WGzQlv9WVhDqWqjVMjFAzK
qYzapCQGB4TBqWOisrXIbzpZIoGpqaFd83MKNwP5+Jp/lmUkizAl7DUXj4LvXAEG
+wduxD1ICe+pErJjdV3i+tfqV6BTn5f/U5hblBflnEB/RbxgC55uYalMHTmU0nKQ
W8kLvxrwUVs4jx04dm9cpWEeQJcFRuxy33kAcTt/shQvkFrUg6EhfMEZVrjnBRZa
iO4Wt3t8j4XERiM/TuWLg4T7nsMOcbu8BfMQU1KKPVInOCELJE6NEXxUtdYSTntl
GFK5/tLrdzwpkEScv1frWPyyqsmfTd2Q+Di1FnkfS6peHBBEMUgze0olkW7nk0lm
tQkX/yFh9ytp0pfigITB5uTj0k+jjh02W4dHMm3Byw5dIm+85+7y0acyKyOq22i3
nMs6ZHw1Z6ylT390+mCwGU3EDNbtvdXpix3TWt3Yu61eoGWXOb2cMUHwNnVQCL/j
Wo8KNm9Qyja8BsrFZgVkEpjGwJLFC74uj2OZvhxfrD+mC1SrZv0iGCE02MDGTdZP
cjNHrgSdxNR5LTrbcGqLWdB8h/XmfEHLD6oLoAo8wKYILgYSk3HjpVDFSv0ZLKY6
Qp4pZUnB5gRr8WiEI2MlyugnLNaPbuaLFfyMylengRkxpaJALaKXgdghpNbmkloM
i3vTfSB5/OG/Q70gzBk5RdoU77jjlY72HAXYydlF9OBAGWkdvhmW+ExMIpS03Syv
MJbgKnMpYBK/py5XZHvjzI2RCEnVZAQPI8WDa3yvVAA6VlPQ2cERX6tnWqgT584/
mdM6aTloXjmPueSXxIT8xHuWqF0OtVQncrcoZIienl7ubMDGN8hxzFnWFe1+FaGR
3KJGt7RyN77l3MNpgy3vRDd+7UwnU3E1VC1dOGIyCYYKn6gvaRiIcW2mIXYNG0wG
aoKj3SjhtSOgofqRH2i59+QCxGraDitW3isSpJDhOZn2kgK+M0kCl6fep66w1z2G
mMvztPA3iH1TW0nfEj7TZHard53gBqzu5lAKdpEungAcKWKlEhd82/FZ2p18L8DC
K+/60QKBPS0hZQCHCSEOD/dKU9s1Awr+5WQYgWCkwNd+ZeXGvfhDOzmumb8WH7w3
RW60e/nWugcjpkaQAp8IUbmIoV59105SRjop8UsGJONmQB79nvNFH4GQjZDVsEvI
rjsKe1kTy8b73Pxj0faKzBMo0WNaltD5HUhuG3IeEajVqjGhblNmFBnqlWUA7EWd
VZ4QcD8ZuQOARqtGd22cjwkK09DD/7EhB+aq7gSTrnOiAFJXQI6n1Ota1g1wpYV4
jx8KBJBoCuXOZay2GSlohm+qD7wCa+szBvFPljcQNgBAgtxFZqWqiZE4XxofNd1g
B5CFPJzmWDD3ziszAohKm4UGGskQ8ZR1V+7SWwM2gGGpzWZTTmk4dgwLL9hzFvOS
hRZGR+20DfmSC9mC/1qiuut2S3pGvw+T4ZmzdTVJ+MxeLGAN9y+deKhjMs9uObSi
k5LkeJkg7VkHcoK8GEzsLfq+nN45FD0LutmfarB3KoKsPBGBWVMWFQbB9/qAvkKB
q3DIzkWlrK5WHfxr20J8sr2er3+/+iV/ezrJNmsqGO88jrblHa5k04HUGql6uIwK
Gwx1yPADJ2+w05dXhTg1JHo+RqleSo7nBXmSqr/Foj2Nrazbw5E/XGnVuRLI/sqk
LL/Ypq1WdS+0qCIpDo6lGXaEpBvYuhX4F52Muc1wwFn7mlwaXWhO8STkMeElIgMR
TKDg/T+BZVrQQT0wr3o9NRjON9yLXUyxnuTrQlltEybJnS+7bV8lwMGvjtM4iqCM
QfWCKsW/MkJNJPqIM8/eF7JqRCfGX6WydHtRrcCk/weFVp6TgmTepiltBrjrmi5Y
sJMMwYoxKjwMaVLu2X85Gz5SGX98AQBmYoa5X16vbvRCPH8IimiHW9m9NZz2BSjk
wHKg+PvwNOXz0POKppC6i2TGs44OdUpX+a2Ah13W2nJxWPIaQ+L1LsgpambV4qHn
D3LQdAIWPKHEn/U2kkTJGgHvFleUZXMf+eoPUuhj3L8JRK8Mc2lhuNouG08sQW/1
2iFax7nKSOCBDFsaOmHK5ifZPAJa7XZsxPKbypPQdIQOA9ttlFCGEHLLxaX1oRyO
uPIhcNT0S8CmhHxjEZYCensXjQrvy4rNybncx1m/PPO5uZF3xOjgSE3HhW4vqe8v
WzdWWyyrKVgBjUdIO2Dm0JLDtAqcVSnZgGt7Tn7rTaVW79wiJaECElU2d2fuzoeM
QvSinorURYPTPH3u+0U97spDN4869dHzt5n0oklD2885ySorI6Mz0oGQS789uRoU
bvKTwx8iwd3U69+qfw7n03kVigfhGBy5mszjePxob4TBD3FtbXHfQj0VC2akk6t9
GLxaiWOgnvCZzaWJOBNRoOoInsbRgR0F/lUIOXijFT30tN2wtxSwAVm2rer7voMF
S+u8DEAfQMIOz0ZZHM9+774RdZ08kbQ6DCAIBIs1kunR3nXtj9vUshVd7BkmcY+e
pX8OD1Msl/AR9NfQKU9R6K/nLN4wHuQLLsphGz+01syjM76OA8taL5pm7feEp4z0
t4GbYWIrAhWYUuj1UZb8LTYvhWRlJTnpa/tL1GEk0BUb/SeQUqHDIYJUf84GPD70
VJMxP54Ipxv0FKQVaI/Xe5yWpw1B4Fs9dGvx7OekpQIyC4xDlE57RJsL38W1ox6V
xgfOXaQJBABx8Y9MUBUAlHiDYl4pUe0FUSESFIA9U7cWxDYMh78kJVd4Ttvqf4bM
0dOfTi6ZqWa5gkuuhOH6Rma6+OTYRi3qNuZDodMRqhmvbNKJbfMjq+sZTvFp0reC
xYV/QYSz1zpP5Oy3uP1o21V3OPV9BrdlFNFhi8VfcVG1GQslaHuMWXmOlukP1XuT
5wwaeGGx20qgTmNG7vBL+XzzHN88B2JTXIjyxYDfvfjpb7Jq96/QQuDLNKrzyVOj
3LKH/prrOSVe6Wnyfqfsrc3X+PiEYBlcBgitTKim7s4jhEV7VGCYU2K90dxVhk0k
ej7obAl+G1uCBtoUUH0M8ICA2EBtBB8Ki/O3u6BP7YjZZAkz3Km3utXC36nI8ek7
URhP9KtaoNcaZDPSgrfQJ5RzLHUGqquT2mDdu8tLNRifNoUtVw34hByavgoxijNB
3uQ07RV10jwYcytv2A2ZpbKoWspyyFB53MBf1Gimyed1QspezWc0FhrtrMX0Gn8l
ToKcy52rWnSR6pSLKD/0YxDfdUg3H+2NMo087qUVS2WZJfCEAe1FbuQ9X1IvHfyy
ANwN9qqYKedkXpzi9SNkC8gdm5I/jBy17vij08M84eXudTiCefCjqMo3uxO0GVYX
fZyoWe49lt+0pXzVqB1Ge4I7WLQFVcSZAoim+28e2MSoEgN1KHGhmqWhT0NR668h
KwICSkAteczupGi9shG/aFjZAyXuoXYN8iRtYKp4xoYk1JIBczsqbay+r6x7LJnr
Gv3LjM92iN030FaBfjIo6jXkEpy34Wj1RdSmy5ZlnpsB/6nOJXfuokdM7ev5koUS
v6qe4YhHIuo6O/dIv9/ujYB3gXYOlX5jocLd6QhViGRtQ6xvWoTC3OKzG7yHZyPr
5YCI4P/C4LqUUm8Bahaj8LA0Oks58t+QADZklbvUXpviht5e99VavEESjkSze+va
ID00EyEN9eSebAyyDg/oxuybGurWqIqPSQyHbZ3+NrNlbriNcUrmZT/w/XXqg8Nb
bbY5IBFoX9lkQFJ+KRxZVo7rECxjcZ+0w57n9h4H6TwO9v+KjaDIgYKOAgUwTFre
aMUyatKGFrQJ+ra3/M+moLcTUSD+Jp29oa2yYJ9NW5lEUasC3OaAm5z+Q8fv+w4T
i0siD1mV6fcL7FDlA5BfPGyZh2LPCR6COwGT/efqnFqeEQ84rgmDp4VbW7SnvwKu
oGnuHuVC4qDTfgsKlWP8dR7rLVVr3/dFVnd8sGJZ0Ov6GxxjxMb+XmaYkoq0VTvv
hgMBQ5LYSX9VoFEoQme9vlPT/gYsLZryUr7+WPqcyUeJwDEGrPMqdbD/O1Aua3I6
3e97uq8DwkVZf3moXcrdrL+wYfLyvy37uEw33h2B/mRZ9A36hhUc0Iz5mkUwjeTZ
sfQUCqm+k9aFRf0ZP+iyive2hvzsHZQrhuHAfX8G00snQJwV4ThRQ++AgoDAW+Qx
NOJVd/FZmRYQCJC/Hu8e+gI7IlXsWfQ7clfdVQxADvl3zBzwuPwbhlzSXUxLk5gs
MkH2pEa7IKigFLvvbUBb4+mvnaFVTHzHgtAzLVGyau0rU5Aq434/og+r+NP+KXH8
3/LZLBr3gOurnIMpoZyb24J8ngQJLuArLF8ZgZhlSegYkOToUvhPRtlxx2uIkOjd
jQHMNXFhh7dhj9bplrmZPhk+NXmyL6MS9TAx0bayy19ojwVmhNqPRIwdi3iUL/+S
aej1Ba8KAW/ZXc4yFR0LYYBUDuI5XF3TIvGQp6/ImEU/M47ajPL+gSzvtnZcZOnW
3UrDz2F7X3WunTCpQMbmX0J5kwR8p41OtptDFHDin1Ui+sZOlJTUFRNDR9esDeyc
+nCB8Wm8u6kOfmISgJSHajJvr8EHjI85a48RMrFJbc8hW3UJnXEPd1TRP73U/HO2
DRCjduoaoldRVM8fiqpu+Pv88e1UymGLIN+B9M+ujOzHYpsjtXsqgzr9YwlTe8Y7
ocy6g4DwpJ0zwe+Ma19t4X1hnIao8RlCZI4X4Qzec36N+tg4/pSwYALzKaRgtsbu
MPpq7GXQg85LRR5trDNZ0nSg0wIiUJlh9UPxqsnIJ5b3O9hPWxa9nqqQnOOzbJrt
vrYf/6KlV5spibdAT/UZgueVmnp9E+pGkqHMpI1TNdFDDy2LerqPIM33pUgXcK0p
PQUlAXkuWM9hDsX+oaN3KLzej4wSnbxu7sGGkc6slJAzEKq4KZpEUXWgH21bQJJS
hADBubrYeCPxWRc9futoOv6k6n53ROcdCpe/s0XcfCHV36F/g5rLqQ39FOCqB4/r
ciUmLKfMwmZPWhF3pTKKZVMBCTKDjYLL5rU+uVg6hJQQl+9pM3NdPCylxU8nrzpR
nhQg8Lb/qwVq7E7+zBPqImqQnBXazeoe2bVHSQNKgNSY8nKq/XlXw8XvNmKt3VdU
z6yr4lu4sgD/zwKMuE/lzKnyU6WbPKC3yuDCxy5TZ++RKbn0OzGzk++E5xoc6PSx
cjYRK1vnYkctVuJjU3SDWRbY3ZUngXs82zSivxDLgkVIEL7W8qLXyI69FwCXeg0B
vSogmmqypJ72dUJNm/1qUUy2rhN3Ys602akOGclMXsaC+Hw53uqxmGfi5a9AqkGT
PsWijrtp3rw3Ci1yaPIenV5xDkSo4Iv5SX+RHw8JtJOXn9HCyHlvfNiofq2C65Hv
xNB5FP8NT+RUsVyU2greexjZiXBe4Lr/M1kNFNDx0P/FL/w61X3wYK1KGp0V+JPd
arQzyGbrX6VdbgFfwcQjiw+RfDPzExmSx079EziKVTGnp0XTUC8K7xxsoD0sMWGf
UvJLEkgdlOkSNFKVWR5AB4MFmHHQfMQTNhZG6Cesd53l75++blxOjbOQEUgtgxqX
uXYwwy8iU++OSNsA128e4ICwa1S0S41mkXoMmh7+NMOvwVHrnAbqMZnGtHk9MN2Y
LhR8JWNTbJcdbfuQHTT4grG6pevRC8SrOcUouG9b2r/Cue3p9FaaVjY91wjUMNO7
WeC9VZ8Ej6ZAD9uax8HBdRioMGZzfDFIWPvEpIqDEoftwMn0WfAHiGIUmo2fQ+Oh
DRU10nTb26XEUAI+UItXHw1lYTy+IvL8WzyCcmofbmy5TqiYaWNfrRJcc47S2Y8I
4+qqEVkqcM9kvxiltiERcH+91vHeX1DMyWY/AzD9tIUI+z0uk7GNHJcZK7L91Vhc
7muuBuHOSvLBqbMvXgyogCKmDQPgCRA+s6vBuZHy13VpCFF/UebCIEWmlU7+GaCY
teB9cysqtFA8xgCJ1XG+jEfPLog5FLBr5H+t+7J6nciiq8Ufaz8vE99kBtRBkZp/
HtW6hxfHd/1lcb7A1zk6Be4NXpDFZS1Z0Md8nvuAuhnU8mW8uE945d6V9VvC3/8C
m1EMMNMi6g6sss+kA17KWX+BdZdgNV53ydQkb+NL7/X3pGfqAUG0NXQnAFkTt/yW
wTNeU/iYqHr9V9Nmz6fm122BhxnstSk+arScrdPpc5kxOBikFdzbVY3D6+cKk7W4
4y/1m0o0qnofbgVHe5zljKVL2UV1BUVutGoRaaNlMiccduuZE2/nCB3G3czmq+wj
AJGgHTqfwb/1vET7AACj3nwCr79/jfXsHtRLcB5QJ7UP8ug328L8OnY9LsoNqUh2
VgKLcQVQUdiLJUl35uZbnbNnvNqPysrzqZwMhagZDgyx6Esur19b9M2FI3mBVbs1
Dfh2BGc85ZJnYc9SjyYwhbePawpTNBOcJtuKYUQ19vQP+TDb4WDTaviUwfXiUdfS
tY/TPDeFxcZzpR6Y+QVOP279aIX1mFzX4bwCblBZ02a02gq/cvvRcL2zgaOCE1Sr
dbHGdabJGzKf5oedLGq/c3D1IYDZym9PhdYo+l7R9vK0p/Nu91gIAhmzp/wcZHj4
6lq5ejQcDgt4dlbaPBSZSuVGmyCIZTyeYQo3Jg+ZzwePnXaalj7aNUdcJt5x2EEP
4yDd80IgqNB0zBs/36e0phwohYmd1Sce5zxuaGCiOXxyurMUFR6e5YqSyq89dT7e
MCCMRFA159lgEbncknvrwVjlIJ1Ep9/pO7fOwtlPO1T7Arlxz4m5ijfV1oARFP0z
CveYxsQGTjhQVkYhzYzX6uY0u35Q9Hc5S3LVHxptXkgvtZOMUviHehnyNjQUl26r
FVSmCus2VQbKt+kENtOBM72MKF83gr0nwYzzOSF4v7RDhdBmiPuwgjq6fAAmqZeZ
WzJW+PJxVM6cEkM3kirD2ODyi95esWvcOaZd713jVL6KD/MZqh6fokkYaPm+REHY
yLS3Tes3nnTyuIWw5zO3TkQ2YFXxNvIl3fEntZVriouotPkJXEZWSuhbdVBH9sBo
xMy7OKFXdSdo7ZDb2w8RQLfCZwSxMvCujkHMtBf2JygOoELi86+fY+ax4GuS1jzT
uimt5vc5zVzCY/L2EQwdxn74FmqkdikZaA9KdY2FadZPPzgXvboeLSPeY2d96gpX
I0PPjHJy8EUaPXGufPTQaB9qZnmg5h75O4f/0qElYQipdLme/XU8S0SF3gxJKS/0
sJJuIuOY3y/8nriBXZf2GxNBdmPhmUHIUAjLNxLl2oHrN34rxAw44CeRcqshhgNA
sM9JSxyNQe/EFaj+oob6eAHt+W/uhdiuAoHXq/tTD/lgnShUFvlLPJaGBHu4cyNj
6SRW39BG3euR0CvQgy+t5SXH8Y8wCKPDmCaDCRVM38RRxIlaYkE45H/iFYkF1/uv
PPOplnnSoLhU6w/EoVRwLTpVXlBviUePKDVxFbOK9quPBDQr9Nsla/atFqByC2Aa
c5fN+yZ1g9o/MrPFWjeSaiWoHNAEhFZpxVrSgg+e3ae+7lNZV+rzAQ7Qgz1Epa7P
+bQymuQvp12DXL7b7VqKVDBsV+YGAMOW0z3SvNI3yOjlcmR59ha3+cB0oZf8zLVu
i123qUW7wQ4/eKPqyIzdky1dhJkMfRzSLg8coM+cBlVh1eIZfXFh9XR56+kVqScg
bFOQXWDul4tG3ic7dXpJdxKjqxYFD9AmFQ3GYYY7Emjm9aFo+tv0eI9S0+RfF8oE
FFxsOtTOJqsYPg67LdaZ8FUMcwCx0nhDYrCdyvNLlTQfOQx32F7DaKG7pbqH4ILp
+15lHDsXpTRh7RYUI0yj2gbtInaj1uJ3M/N9Exp19cgMxMJiJmSeP6Owk3Wfy+gn
Bj0aMpNgHBwvoxe9kRW3QnWte6QHE1Zx0jqsACzCexmZZ23ynXD6jaFqEzIagtTo
Xk3W7INbYzXsTFY4X7tnBS1Ubmj8UzeFzF6aWWNZRhCxpJzMvGoPPMrYlw9ftB9h
QV+WNx0xGYmrin+M0ng9Jirt5c+3ESJJWL0Qwry6L8+6WbZx99BuUwnpmeEyoLXg
Xy7kboQeNUo5RuBY0SMgPsB0WEB8jxETyuuXNnPq95lOIP9M1tblJ7YRtLAD8+N/
/qWr0058BwjYsdxvcHveX0WZtglFu7BJ4LU8re5jEc2tRHdM6TJ3TfCKPu1Kpzxz
Xjr/OSXwRtxXtddy7+eIfktX74Liaiq0JIdMWBfIjkb0XVDkdqzneXHlzmKAQiyC
OW0xVMtHq5MPNB5BVfF8gNatMLTbIbWW+3BACVj2/wPCLfvoDBRK9KdxmJpn2iDW
4iQ9S7TGJeTm3HDqu+ZCSREvhEyNb9j8778tOBGrkMdJ4Y0blKyVTdkcLzsSV3xp
PgBPXKyTvgR9fzUk+I6obHPqWYDjB4+/ogzIPEzDLVlrWf9TIXVUQl3ad9Va0mNB
hiFryaiw++D/do4/RlJZf2xFR6mZvRnEAO6X46ieVwC8yTSd9/yit6pFqCtZq9HT
O816pxFSgchTHjAUNSSr7CXtbgM4Kyzo7Yzcwoc/PZ+7Nb6fxCmY3n7GDPyK7Pai
NeTnEo8ly7nhrU6ZIhZK7WUNNqrcsvixuH1zcAW3RdCZaAXGIS36zB4s1jELn1XM
94ZCStB/4wWIRJsrpWJGfWJtjs5Se2Mw6WK6fG334c7U7228vDigz+D41HRCI989
cFD85xx/VeltqQ73L/BOxcu2079gad8i5+2ilGxkicc4Zkcx8bqUc8nIpS5mnvav
NYJ7koXz5L5FLAadTRuH9NsjOXivSPPj4anhzilH6SvxdrPLFvgmqvQ/mBzpRdVe
LCHphoxRrsNcbun8WMCQncZ5hSTqhNWzc7Jy8rE9Ai7hRlCs2+3EU9PN87pmHz61
gwgqwbus0rAXPCQtucYDBj8quTtrTwQIP73J48HQ8AZV5RBoQYyCWvGGWFj5mND1
eYOITgqRA0bCR8rs05VxebnH2MNFmFdHZoL5pf6wFfPYt5a43R6Kd1GXYwPclBJq
YPwk25fZWEnZCNinXkz7FeHyuDUi8eVqzSYVigMz71BicUmDI8jFZtNdRhbOXDJI
RYqmzFZ/1BTd7/EBkSMvC/oMyy7G1mRBbZGGuOIiI4ZC1rfH7E9mpaNHLMbJqJD4
oC6tAWq90Fenz89xL3xNt9IDgUn89S3zY40oN97r8p95ndLcK7sMCW9p/WGorOyN
5Eh8rmapdZMV8qDAPUk9eJnMtDFtNryZSMdrb3sYhAzPFCzJpdyf6mHr6YsGSFtq
5kEt7S113PhvNR7kVi+NtvuGmYFsgZKficGOKI0XiR3Bl2cluboKda9/kF0gLW67
DQXpWLpzWNNnlWNrBYKHBCrCGLG97gMCEhtsYCiRkSD5W5NPTdMEZO+KMfZF9vfD
OquMXjHZoQOCS/XijYlYVaB+Z6ieB0ODgfN0OlmrfLKPf9aFavoQBJoTVM9NRu4u
FDS8NMDOgM7xI/5OC/2hNZ0xiFan5tkHQgTiz+PUl+in+w+FJW4CpjLEkZh3/5sy
5X+iGdL2GjKnbe73bsywDZEiTMCQZyMTORoFrPhfan92LfXuLr7+umSLFtuAltFy
yk8Vh0c3WNXXf/OaXZIoU03QnFVyxTls8xF3WZgIzmga/Twg9J+qiztw3Kttjgaz
er5Ml22TmQShLk9tZrA6SLcuKbgi9lwMI1+acUQ7JPli/rB11C5avyzCJyB/57v2
z5X85CyuEzpOaVDpch+bFfg8NOMQXsWCZ6jYy7L9qRAS02H+TnMqaY5R0RZU8xA0
Go0X86XSXwud5Ec2SYVzYnkA8+EJPWeuyl0G8DfcQq0jP7lHNdUcTnPGnOLGNB2A
yiv/C+ahcT71xo2Z2OaJFDARxiA9bMntGSlriEv8Z21FZ3O8NYYFZbybp7zjaaWZ
qvKp6jOn/PrEeXiP1n02s0kZRuQKFV9+VXHf2Xe6eZqRmvULRUreV5S10MOdI4dH
Z2CHLFyr2BNlppEskL/2tJWpfo5kQNlKZOy5lDt2UxUaTAcwYUN8b9cLqKFy+5PI
XQhdxLtUebFCqUKr9enta5/hId5wd49kjItYHoFzls0c484HX0S7Lhf2/ZVIhDYA
XLErco3SGNeCJdUouC/rNnKUPlf7eOXl2EgKm63ZJ2+RlJtjsOqoNjHed0I/y6Q0
TKcnJ1+ZpzdouJbWmc8HJDvsKEwzBpyfubbunMuQvM/W9u6enOsXbNw3oTKzxi2a
enJFofEk1uB0ZNVA1RLIFzn9XJlwXo912hik1inQcO6b4d7Vrku01vUKqhZu3TAA
CufS8CNi8zieo9t9tihuMuwrzDOS5Nbr++si0lI9b3EaLB2I1T2/aXu+GVdj5xPd
T6UnoSI6qcX14wKN5ETh5LT2qN3tO28wyojtGslN18lXBkTDVSp0lv4u2pe//FeL
8JHKhyDEymgJp6vE7FEUFrqj8tHtx/49kiQycVzzOFCb8/5VvXsFocNI/CuMycLd
QX/BYwIzZeOmUf+ouBwL9jT7dXl7q3zgrF4i+GVhkHyBKmAbwXGrhjXM1+7r/m/R
d0X0k7V6mwXDOm3QY2JXDC8+cJ01O+f0l94wM2xS8l4CKB2DYlEOT9zkkyWt48rC
SUML0SGluYROQSaKJ8GBAj57a5pooDnpbVGkfdTtNKAZX0SqGIsbdVc0FovVETB0
IurmOnkqc8Uczh+KE2xPpCeTX119xVSiEL0PHF261Z0zClUihMsHWbHfTSK/Aibg
7SK3qJvLmyITI8BZ0Ho6C0+XuzuQ2MTWOKtN0/ypnL8V7xUtYXoFWd1Zc62nfb9O
uJUh7I/ynI7tks8PJY+FN8EoQ/aOgkFlb4nkZ4KWud3lpGTe6VQ73Ese+geBCYVV
9quGVoi7q4kfvhk9JV+JyUNCJQqfOQEbHiURoJme23PvhhQVrWyjmI1+Iza0skhV
+bOaICnmzWm6aw5wH7m+YcYHiYyhgISo4GBgy/FRHbagqBOIQt66TjuyDpAwtw1X
Iwu2eJabIETdG0of3iDZnVCLoztj0cvEaUPozKqOnJBF4cMQiGoJvqtgq4cLPDwv
cMigADzzq1kR4nUsFAX0N19Dx3YxSRDpT+9xSGRKXmtAokodifNvQ/1NqlOqX3Y7
tczdv0cOK6Yg47bKmDkBuO30L8bT0GthGGOINd4j2Dj2vTobCxlLudWY4uP4LSiF
G/EcjGTftGzmCvrY/GHd5/ivLL/7p1QtvLxsDcN4AVQH44OuApI7sAEfY6odSqJF
iL/Q66RfSuepcxlbj0xy/yxD0V2L73jMXfnSNQ1j8gtOZV2e25mZhbkmawCNfdxJ
weLKvu91NAG/nQP/QGuuxY1tYpcnrZp20Hs3txdg4czQGL00oWkJ7LaiQQdAylWy
hOi1wxGncTjKqnxQd4XOxN8r/v7oEulrVnhKKe15+jby6KB468pt2WxpTa3Y4nRi
EZLeUovxjZCrgdWOj9v/c8N4+j35+gVgYI9HH3VUJsVmcwbrfmBYdx3fb984PUFY
btu014z8t/lsfeNI/pjVnXY6caWhfOe9G9ciMyrkY32sIdVDNCQMgtq5wFHGRSPv
Uln+5Yr8tJwIMpMTQsujidQ4lj9BrJeYr1MBCRGJJyhDNZdGqHPVxrc73wScc3ec
lM5FaeiZin68dEMZMpH0Uk0BBJ3xLuGP1F/z+XL/kgDU2t0arqKxIh8GnsGoKPRC
40Z1cuwefyFxRoQsPnwwvHLQVv4M4hgIL62+vYpwtdizOIGVy73vyi3VA0iLA7BN
mwb8mKiBjAK7Sh4ECQMKk+3okaNm7fUFBzFXfFL4kpVwqPU/69drkz/IY/iZvIAw
sjUI0zfSL8JENoIEwoikPPsxbeLxwfmDul8XChgCjuqWt7T/kP6+9nc4nAXQiprp
MorW4emccozcsIyuwIwHh7uuJBeBfjJvfzyIFshaWKYNs9jmMPT3NTMXvxpT3V2X
eoDb0PanDFHi1jNSZeTv62xi2Fsb7BXj/i9RYGRH+9BSV4yD1g9+gkrjfhz6NI/S
1Rm89PuE4U5l1HzIzx0G6X8/R/BOSXEJWxhQi6MSID8NNRRoeNBufGmzVAG9qN5m
+0QWhpffmeXHorJWtVZAPCVgnLgeWfSBUwDCIk9XPXl48SaF9jskDs/kFheO8UVA
GKa6ihaJcHumOuZv3XLNVhsMiZtSwQ/yzC+6BI2EFsmHBdAqCmTCUmq9xzWPZLjR
Pws0clyoL4dsdZqwK9Hp4rjQhw+5vbEh5Pw+PEz97Bhv7F9lIlenOKpNdzpzotdr
VaIU4Z3xFNKSA2f1E8PDHN0nLPiUmmOdNU2RSW61a3OmVrpu9iBNANjf+SxmwV1A
Bs8WuFlJcsWqPiDq8zKAcsI9f5gxZxj5lDIE2Kl6PkZJL6NSmU5sVpMaEvrdXJLu
XzBvCMPtQz7WZFpQLIOBYAtlPIPKC8TDknANjcHbbAxk67ofAWlxsEiBlNb9I+zL
/JIF9rMmZHZxyMycPWev/IyMMo8eWHsUxKFa1q8Nx6CSmU5QQcieK7WDbEymd2K5
HBR7Vmw3EJFAoc8DQ5oRircF4WqAZtqDNxXTQgPcqdrylYcrDSRx9X4PMYglMsgG
RnAp3f8vbg7eBhBAj7T0n4RXCyaHlXMyAEdGC/Q2EIPUMIHIqZGvrHc79Z192OIQ
bI7Avv7zqbM6bHrV4ESa1ez/FSKdgIHhFKpDwibbdCGO1ZIaKEnK66xiA/zn5nUE
0OSul/4lcOXk8sI4L+i1MO5l6cx7q5BFIydZxhF3RLcxW5MESg6JjqhCsKVMUY00
lu8kLAXTJEGJCJ2D7fypbKuo94XaR5jwbw4pqCGgHdxSYe7UJQSeMGS9kcPyVX7D
c0/YZqEW6grxboOZUoQynkXmCtF/jkkAPnOLMFZAOrlYICw+3s+Ziqtupf+SYb4A
vDe/Y5t9AHLBaFEXH4KfkMlm2P50N20DrSns8VEGP0nyJi3l9EmSX2a/OElx3Mnu
srW8CMKj/MlS/vUJdDM49vubw1+0CvEs2v5Ks5Wcrdkl4APvc7O0IspbLmT9xIvR
EgHBTe4XBOyUd5ZduMkkXbriEGnvgOysH0lqHVUy0R9VHXAXxwpC+/W11lRbK7+4
GIgs0dWFSZw0B80PBPnQUOEOGRIdZ+mCYINwtgnNPMiN/HyfZHBNXacHVTVlbzb4
tilbabGETAP+rdFnmYtj66TySuIksNRggbzJI/ikERQrt1OabCeun1XGAMGku37E
61H+40+mcPnktxL+DgjtnnxPac+YzUbLqFiNRYmiR32O5sEFFutRNrfc9wSO2I43
KEJalpE7BC0p5AdbRxt2cneimg/BT6vUcRo6DVcQrp3SCqngz3Qv+1+ij5kNaLPl
Exo014nCJllIOTr0C61fr46ThiStFPSvVd3IHdMoEb2vUBmK8BzKryJY9YIa6ou0
ksuLzBIjRBi9GV5L3juCKOAoatqlJIuJkasBYqSS0Hba6eXUPN4othsvp3nnHM+n
3ByehUlbhZXeEojyXXX8KozkUO/N90ieFkWBmXA1Tho=
`pragma protect end_protected
