// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hsl1aB9bdZmnx20wPqLuoKdRFNieV4c/TRDYvRi+YhS8X+e0U2LQdRnYCI9QOVze
LygwOdeDL9/MVeF+gawdKwaWpw5gfue7h/W+Lv+FbEO4wosfHMZPb4VdL4yNxgmH
xUwl3Yz2yFPAIyN80Sx1t3hMFethwJ7qopkCigQ/z0E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3360)
6oMwxiT0qyS5K9FYDHR5JMfC/zdmpfcNmSscapC1hD7g+wZ4X60XsKkGSqSwIXXE
dDqCVZYtX9nqxNtFnMMniHnm3zJT7IhQK5fQhJmaZAuqGm4dqDtT6Vjacx2bne92
AqDmbVwF1rJ8Z/+yzGwh/cBnqV13ntH49XTlmgDt0BYCgIrZXWjNymWelundAmhV
m+mipLtuqS/ooW4jbknYR0Tyrh2psuD+LhNLSDLxPbEOkxFKY8RWWQvIdvk1FRNb
VgEjxm/0IUCBS/v423zJgTYaepJAhiz+GCBkxUXzh3kSNGdlh/4acCkp5ZV4JpOZ
ybO1TN1Cwox1N/dQQ+eSFALiIAnkSZx9HZGORkCEWwWgZ+xkf/e/pVx8EkdKig/W
tIpQMWTQDiVgEcL4+n46gw9XEjplObuxM6yMqcjWTfep8et+toi4sIN+Zvo78tul
QRJJzsydQYQR5n03HaqtgQ69uGMsqNKGhiE0VBoqWMNgZHmuZV9zOInkSZmcasqn
V9LpUuICt8wnVTldAyQhlqCsvjluv5GIHdwRp2/ArUVklXSrVTzkVyhMRGmyK/av
c0E1aU3VWEJ6U70DPcqj3U2If2pWY16PsrrWdCM1tG5qJxPYN/hFVXQUVvVc6Ikn
mFWgPZAybM3P8Q6BWJs/ssw6S4gs/okmmi5nQRiKo4fywTolZqreMRqgTqCy0OYA
iuqAEvFJ76otlPby0vcUaGTg1sz1FIDJWNFze0Memr6jQsXFWpevKf8LmDmq+GCZ
VbubDXPtRRTrZB0YrcgBWNvT/dcaZA7g5xaDHUzudmzvNuTwsNZ+CkwTvdAMfsIZ
72u1QYiDcqPk5q/WSCK3HCMCqPKK27kjx0CDRtt7xkl5k4IRgXfNgcVDsFdsnrR/
8wgPy+JCGZQdTdFHX9OezWXkiHHiHAN9DepFUTLJhK7L791XTDeHwzlJ4GwMvIDE
wrT40PQEMMfsaSBiC7Dcfq/0zHUGO0WZIpD7KWwkDk+62Ti3osC6Kl1WkTG2Ollg
y2LMR0iInnBbHoJh1GHtsQ3M6WSNni9IdNtGrT32f72fVWcrfm1KBQy/Jbi5dC8M
6b/F0IV+f2lotDXFJNNv0CP+ntUR6KWM8DdAABnQUxlAv6vaFki1EntyoLdmd8S0
e5iLMfAJd0MJYLVGzcMSu2Ze5j+kxdi43XvC5ln51kdXcG64YwsOSKYoVts0I53l
xqLW3+cJCKlx5eGEyTOsEneOjFgVTRpRPRmD+34EX9Q1tq9ZbzBHFhXlId/cylop
6dDmUpAdIrQTpAG1Pp9sEiG7QrudHv/voeA4wNY4NU+z+Qzc/lpRXqse2kQ3L2O1
lfNzAO/ysZ8Vu/U7XGdRn1foT6vrbe2u65Qe76Pkhgekil73L7rjAPmn2KvYVHY4
J+IlaJAnE69czudqSa1ZQ3/J5VLVBs5Jr0WXQMQuN8T3IGDbaL00pDe7MNQPc/uK
vzhO6id8yRAckfISJo7l0gK7M1IbO0nVPQ4dV+3T7YcEoC8igq9OB776J4do9+SU
uDT9OA28kjif9WDCqNBoV7O8CaiMRJ8RmNNFjd5MS+8We4OW7ECun6Q1ktP6W3hn
hlt9leRoxEFhzGo7qjG9UohAkHd43YLdDWa0qgvscATqpA3G0Docm/NbuFX0WKuc
s3cEG/IQGekhWSW0k0OR9AyCi/B4YCRZ78gxbAvkHU/x7YHIU6xMx+YWd5M64e/8
sK2l7R5J/pIssAljYg0t+456OgHbh1yDrnRzC2Uv/11e6hGRduzrFlqjKCJ6pP+o
423eK6zIbtNd8CpHjzRd/1K2eAJoMi95E2vWA2QHm7QLb+nmjJx0dpIy0SCchDTw
HcudJGE+P0frbgeVVKQ/G1riDgofxO/rk0W1P2i95LcMUfPLks5Jl1qtQh8cJBKl
tPsBmm+jDwtaW58ZAIxy3hVgg4p5Zc2ObHBJ2DWcg91vtZer8OVOoty9GBJwMvqf
KWhWqJO38M8iBJZ8LlUvN2Qc73p8vCDWnh5mZjVzLsxuQC5sFwJBFGIcvWqqCErr
KyFYcwHAxp1y3yVIBSk62MV3wSwW6ydkcs8cMIM2+55qFnec9ONS2DVs4MPPTcW5
FgAM3CLgC/sxjSLFqkS8WORWhlnxpsnX/1i87aY9DeowgBdvJdvc9a4kbGtzOM6c
Tv+clXWhfrha4QL0ByMceU5LbxxfAddzp+KnxZ/zNfUC5jgLXDj7pgDdtqncbgwv
HKAzsudbCCeJbT2usbhUgTEGjPaCFMUAu69oA92fG3Kal4Z9Xt0F99Gryic5R4ly
iVgIDRtHUsPknhImfsaetu9N4avQMe8HVM43LEBaylOJlGXnv5gGZt3izTDM/rvZ
S0yKKMAW1Q03OdhSGWsoB3a/CIVlU973mjdBynnjlyL8Jv//YefdBi1gm2mmxgcr
hh9BjAXA36S8zUvA311I2J+2y2A+eS5PcGxLfo75nL159oHokZkIX1Nc7XDneKdN
m3dV/5caLkQYyUhx5inugDVN/HcL78I6xjpRkplObUuXdvdQgYF3J601m1Qio+sc
lt9O7pd+diEynuRK782TNdT3928i4jWsuoP/N1Q98u5xggAy0gkkYmYpolTo7bBs
FmQa00PtT1ZBmPQ4kzVW81pPerVW1sIxOxgRKovZE4ofEtW0LPXwXIR7INHCg4mV
mEwj0br4F4Z2X+q5T0sZE5ttiR6uL44o9UzIcX17f5knr2LV/COk1MDHdM9lP+5Z
DdkIAJ6CUEqR5dbsrUTI/kigsZ7Zlz5Ri9IYGXbqaXEPBtlcTTjA7ppqE3Qpz/px
vifA+GloVciXAD3eqGRrcuZ/ilB/kzputIUtmtqN0zDp3vfK8dz6GV7Pkqzj8pco
3s5xbuRfb+oWc7qA+9INRciE10WJ0ymDccURrYIfeCLs8G9y9uUY3pzgTey7ggYe
ybhYpK+xOfKXLLf7VNlJijMPgF2ox/x2YIZiHf33qbm5UaqThhSDhwxLLHRMZ5mA
bZv5r15Hr8KN/cpQl1MF2ZIXRJ6lNMx+4xkwjPUjI/1p42oLnCx49/rryNqgdzSV
nGfwPoxRwF+lRIMJMbmjQglTtlt/XsahzqWFHyiQJ2PVJ5Sg3nAhnztW9o74TTbM
zkw6Ef3VSlXUWus3t60NfJo0t+iu4Y+ycFW16zRjUJj/THjsNTTDZB0DpOAwyw1q
5aKGuJ/pCUeY0vE8YQJjfet4a6Tfi+SXJ0400zGTtELiajGKwZ9ZCZx8bWR2n9xZ
GmbqfOci1w9KEy2hQo5K+wlD6ZOugzgX/NW6cHDvtWLrF6VELeE/cnOzhXiO6PFZ
WR/uVS6Sbw5S3QVHo0KSnc337uTYwazWk8eN7fqo4Pk3T3YZ4EYa5dzUmwe4XRa1
Jc7LKQg0bsvg1ULcKsEPxFAtXs1rwhsCYGHwq88USN4wpIq2FkpYSBZS4KbZDNmD
LmLZYh1vtnb6qpCjUXi/U+5IpuNmN9ZsHTckSx22ksq1QCDzSwyXKsf0zuBAeO6e
67JxwQPTMxmYNepelVP7H7vH3fd2lPOulnckWMWDeou8TwFnw4+hJ5NvcJhPoDlO
YRGXCVlFiotEdrkHBgaRn/NS4sxHnnVNL42RzSE0c+QMfW1YKFKNsuclhcEYQ7EI
x50JaokCAUTpG67ixuBQO9raBQDHg5tGDWW6S1/1GAf4k05S/0SEaYVVwfuTp1Vl
ywdAbuLjWHl8H0mSVsT+Oa+OaVdcTlqLrtwaj5kLYPsVJNt4O1ADHbPavbTKe2TE
kw4NnLCGbZA7/eRq1M9hxZr4G9aRP7baNEAGLhyFZdWEWUaV3AQ2fVz3gAi2bnnu
yunR0Wqq6XIb4FkniLFHku0FHYWGzLex1EyJG6zWEd0UYo+4w3bLjeQlFWaPt2pS
JJsZnWmbfM+3VR0xejhOje3nV3VGX0H4cJTbZ9MJKjGlTH+jGm7YPPPmUMeE7mvF
ASM+U4f4tt3v3rNxb12Wla6af3vST8eSXPHESrihx1o4ggkZDn+G6GIyGS+9Sn/O
YLSVHOI8BfrwKWg9RsczIO8543DOg5hUvaJLjQj0tRfBufD8pvA+v0z9VWpOVLNQ
UdVEApXWtql9LD6ttFtT3IXj/sgOd6UsLCwQQcMFog6DKdZNPvaZXtYBYFJMhEmM
bWOdwuXLDF0A9J9m10RxoNsuJ5SLNl/kFMU9MRi2IhTBcZdsCXfZaklSpo03a/Zz
OHnFLPXceije46QY64qx4LO4SxSa9Eibr5w6iL4neDgG+ZQg7K7NqhJxTHImSRNG
RZG8D8wfYFol2GIivvhT6eReNxUX8AJ/2vztHX6NHa08+A0kMLuwWgL6C8ySkgOK
kxsrFf9s+d6ALF/8phXZQAPCyUR6pNK2W7nxQgTaJ8hTKMFoFaHO8YZqFlsz8IDg
QvX8qMPYm5rDMuXPJgKetpV2BQ+8xu/QIPoVH94PPr5xouSHu3Q4nT+CeTkWx+np
`pragma protect end_protected
