// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Fc3iAEH6XKl6MJTrWsEGHcIzyOno6afULPreV+AI/8x0XinyYHY8/ywYWN9P7Plq
fugZ3IMRi/XX/EntDNg+UlrCdQnLcFsGkDsMGr9/jAvNBUrHn2xg3M/womoTaKTt
L0u2uE+Oyta9QQ3FCxMyh4MH+B1OCDppoF1mX9fvfBQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21808)
agR3xcwBqc6lCFFdKloZKS4Bh5bcH8fc15UPnS9+g5XBww91CV303A0qYCtwQGV8
6C806lXbWoy7T58s61U5D8eExayusAqf2M347rL5aYGsTe97Rp+K6Pf1xVWfAzgO
fUvNMU0M28CaGLTgosj5al52JSjyemZyr4+g4e/2bUEsQOFWgnk6lIsAMiAIDqBm
l2rHOLsvfbDK+K5FbLy/FhwwXaPIjtOssmXmZ4ces1t00mc+hRWR495RDu0tpJNm
JGQWQAu8EmO1KSSpY4ejLUmGBEHIw05Op6I5AYnegviwOc36u2meOzpGvfBqIalT
jgXDais1y4lMvQ87tbDVGR1O8sXAupr5tbnEhEb68sK43Cf8d5vrsVETD/h3wJUM
jwiAQcUmYkugL8FAESNQOcFEIayOQp0dbGsLjgzqu4iN6EH3iEZgieVzgieNcIcg
jsK3SW6b5edkuyh52Ggx3HKGGaBFiDK67mXAAbgPB0jSE+N3Pv+HMbolagUcGt0m
eVywFJhANfkmCsxL9zIVsa6GzwVeQ0YLdmmHlrcrDPOY0/fhtX+eF3GbXCTwCika
kDMO0ppR6nS0N9zkxhP4DIGJ7HVMxxeIsRTy57mVFN4QVJWf2zNu12hSKUJzYTDO
qka1P+UjlqKWKGNk+gULytfP4DkvPVs9gxFYnJN9CUngsgglDnI+PpnBjdoNly1H
vJzdNC1YyBFHVGiFTojJBsYDOGoFYyTkmxmFqS7qqR2SaeUCNVRx3SM0Oe24uM+2
DK2J0mUW7H1wJexNrzgtu7IAunJKR2THZqWfU3TvQ5G0tH387aPJtGVIpPMTnyxp
sq/atHd3PJB+uIK2ec5RnbOJ76MuAyRHqLYfvNbLGRbwuI+OxdtcbI8q/Qr0T1Bb
3FwtG2gEJPUxuM8qbU7LKupYatts3Z8jO6BhCgcbu76flT0Tb0bYICYHBX84OSsk
EQZFrzM1jBukh9OdLSF3i++wNp5lHQo/vvFvU7p4BVY1xK+kadTfoJACuyuNNylm
O7E/vU+Rx8y4KvD/KaejsGSlX9m5zlERYJ8cMEzEV9XGSa5tUj8H99h1vx+jO5Us
BIWVYnX3ZhsT/4ttzf7x1waR8VG0rX3746AmAobRMHzukINqtEwt65IMw2ZylZrF
+2CWOrbc9Hu65fV4QMXgjC5reKCacgRrNJkM1laPbik4lxscTsMuqq2Cd55Hgr0I
BngPPzQhCYyRDqtqE6j3en28B7Bw6skWbaoF1M0vJaXEj7ND3s0FhYsQ0V0/Yn2u
7FEt7AaYEpCuA5Rgt8VGXW5PMwrjEvgVyWiEVHo8QXb9zezN+Wy/Xp/TKFkUiLug
x5YyOoXwVuJ6kyBigZbsIwYOwf1FsFBWl0YZZraC2BamVdMnx0CwuzWQrqGunr5K
Q/RvUJUOyIMxz9u3ywW/z8O0tm/mTIiGbcPsO6WvZpAzj9norJqi1yvqHfECq91m
5M9xfXZ+lcwSyi/3HZWBUmPaYujBWH8lwOhW8bi61Jjye9YNSL2e3t83R6S9Zb52
LM/kaEfbgoTPomB3oHhSfn+xDm1yHhIdeTOkO2GGhn1ODkmG5jo+r7GalrwcoeVG
OKaxKlLDFBxHz+fOn7eCBTnIRNem3xGSuzsyEIRwLw/dEA6/vnhA1+1BeV7bn1mw
pyvXkH6kHbfUgA/06oVA81o4B3WoLZfFxWQN9rTpt6v6pBGc4XM9MI1gbYxp4Hk4
whaL6bqh7575/w+Ozxon7njakfItuGqpdjg1Z6YAX0pztXb8fsO83FFmNNc0OZUP
NIZ/NIHyx52SkS8T2/p5vgK2+hbhySjtZ/yGwaoRsepFpLXY0K/Ti5v9snvmKm4S
zrlbqmURk9p7Lvb1HEt7Ch0lKqRn6scBPulkcvNYy81+uWBcB7xPVZprFeTrMJU2
cETV5ENK4ETqsOkOL7nlW7siXRsRn30UYiBUmnp3dXkT5pRI0F/sNGpLY6uFgM/o
f0aSaBVYwFh4gU231XeA80C8WAVdOK25rQZJLCvfT4sBSQcyH61uxfnW4rJBJFv3
3x1gTeoM9yDhdxxtyFhFxF5eJlxHBjrorn6fcaNITs8LNlbgXYfk7D/prT/0Yy1O
2ZNM47qKm663gvrOtj5WRkTeIoSyk2knfLS3XGueUkDcOHUIKU88jc7CBT71kEVo
WxtTiyHIFoypr/+pxMR3MDIY64J8zr2y8fZ+FgQXtewSOpNgYLyTJgfCmxUWuZq2
iXIG1EBp9C7O8b6pLXf0GV62Q+CSS4tptZTHXu9a7Z9pqK+Lu0IgoWwOIp3PSe0u
ueVtzXG2gMvpbCqFvBa05jH9OMvvnvnP2a3V2Bp0g5L1l0KPOYWoySJzog1xt3lu
n25uEZ6lWs1svXMthz3VmohNog0dP7enHQEOHNPXl+oDH1i+f1hoDoMOMiEhf8s2
BRdRePITO1qqyeAUn9vyVAfnOo+BY8CepVu7CcIglApNzDhKNiirW6NjFo7FrV/4
zsKxQaWy4RfP/hUF8RS+YQ5LnxLX6IIYwffbUDDiAlBWNEr8fCTgVH31GjOdjZo6
kq2NSy4o9TTaP2nwpydduAzr7UjpFaMSr/mpSzeo4TY6F5BU+RSQ+tCAr7lH21m0
ESkgbztuY5D8qQXJ4GCMZCPKlhbAUVuXTH3jdjX7TPhAlc778cBisMrRmRxsOJOm
N7JSj0/a//WuK728aliaKaxqnSnvgI2FEqDr7R/jo85UpFKBibMZP8jypTOHArTc
J9ynphqsIn7YdOBoiqHoR0tmoAzL68uWzLKlfM4dxS1IHFnUEkv+wijwV47ISPgm
DeFTurXPkQWIcCg0FJqJB79bE/FGqfN/EKmVoVkiEdzMZjjolkiFF5oWWLvsSnPP
3lC9UFo4KKp+NSfUvDH/qMhC2fiORF11RJ0vqzVaWvWcTSTOPq8LeZIguEQ9vwj8
Ivba0nikvLBJYRGuxGSR4Xm70/eoVsiRTPQOSsucQmLxKpMrOJs+9kULPSnrNV0w
/+guFvxI1ILBCwW/xzIoTD+U0mJfNNjjw4d61bd2V8P/MtOU1tHQ/LZsNovDLDK9
TwXszuKPpa8iTNESDn4EWFdPbY/nhhc1dIp7+TS2klqWjabl69BZr8qqnclj7b7P
QmFBx9i/BV8Cfm1EjlH7HA128Vj5+O8iy+aSBhc28QOnCXWSPGG3UfEYHvLT4wQi
+AILrWhUwOKy5LJlU+qE8w+BsSSrhuN3yCl70E4vZieVs2LoPAQGLs3VFzrpWzI+
gXoGaUcVGKiUMkO81SUOZAAvuZ16/FejrAYeWMXGdH3uIIKynb2lFX4UilpCv/lk
6y/ZTn4E4fGM8YWdHl8AevqvofdkTsnS7R3HuIQ+FTNP80AIF6nEi2XHkJR4fdYu
aiZxJvvsUgZ6qLzeEMOG3WZrk24PUxc1Y4AUNnKJcxsgiUMX+jfpGtXMVliAVwif
en1iQeROal4zjU6Yayo++oX4A4CgpExOBlS/gxr/H9h09bT1W/8Yx5R+9MMAXsc6
cNPsvNGFAnES7w/cGI1OaHeID0qqiGRD68Bla72CUxAoKggMoIJv5skj6AhumGRV
6s34st2HFXQTKFCr2IfeywSfd7g4tq93W1oibr7N/5Spg0nggDsk6zt1mdgBP2Q7
bkPMsc4PgexOowqIyGE7F8oIDo0/POQ1RBTXc+2aRb9u/vWSFGKMAwGTl4/WTE2j
FaX0usbvO0CwL1GgFlvDpcMxRX7v9vWe2ajvGOhlavFUyiwsF9NObEmDvzmKitvr
D/OXCBM2QSZS7h49ZSOB/x4dinxrMbzkgGycdu4oGrC4npA3F5EbH7E/qU4Ra+iS
4LVw/D0KdU1R8jKscVH0E9DyjDeQomspM9H08knJgtLwJSCCwhSaN8CpVFjNExhi
65JXs97zBjNFcoh5vA/Uox8wtciW3VTo13qsaVVZKZ4EYGfIx1xVYR9sTJG55fgC
n2Oint8/aFn/XFyFL08wBe6lbaSCq3dDzeAsgzuYxVaPgSOCrk7x3896pYuXxHtP
UJ4xOtrPWMtICIi2yXvBDO0JZFda1mhySslOXAF9P/xkA8Wx00R00ebiyBhlBSXe
Ku2m+fm7hPJxmSV+UJqBQIqTd3T2eAw7OyC0XgR6VgmZwXomW5pjmtNvdRBUj3ET
DyDgxnL7V0oj+7FrjhTJU/yfLUcn/rE23kKS9oYzytfhSVCjomHejpXow2hSXuBG
Oh0pHzkxbOqIu0E6AQWpCjJ4Q5WsVRWffnyrCmVNSz0jQuwkuQtJsatp/5P2Zg5Z
uFRpnav0NYvsFmzOmj92hI0H8JIshxeBieZtLdcypGBdiiLjXZGY8cxNhr1T+Gga
XBGGAb6SzjplloarVWO9ihFQil9sqll/H/GuAurXpLYnu2XCGaMts0NSnre6hk7G
01Spk0DVOpCL8rSV4ACIa0nr2X/bfJnthodlMfxF+M0Zc9AcjqjzA+VwZiw13e8L
n+1gjNtjzHiZDg22jdIOYibY2pOxzSrgg95X1BFXfa1Hnqh6MTibyf3sNtcpVXfP
56tGPfg98Z7sgRMJWxbS+lSjF/Fm6mLiaw2WFGUB4ZImgKHgmoKF8GX2KEPQW+Uj
tCzJWm4IBpP2N6g702+KvVcwb5ufqVa8UBnCPaW5E2IEHCg1imXHo/TRHVB9xHRw
xaY5C2Z/gEVuT/Fq5S1GiEV+0jrZZZcfaOf8YjL+wGzC3uGoXeBD5Pc/SlFuecXP
+UxVo/Kbz2Kr41Hony25MMulOrRdUedwV6/+om3xmDd8UB5rrJNVlhSKUPsH6n4n
1lDukmvqZDvzS1iT2R9qhldlcx4TJnA8G/YkrrRh2WynCaDBdwEj6tDu2Z6CJQfm
jgEMX1orw45vh6WNu5XIIb5iEnUg1fi8J1r+27V8QgEyhchDunCN0NiyYRU9mYQa
hWXa2nsv+w5rO0UgcXr/U0E2hI3NzvUa3cf3ViKlDDCVu59t1QZHG/OgXiml8y69
syv51HiXvCZbRQrSE6j2lZdMaQWByAkxJG5/Xh9KsIUux7j37ZSF8kpeUCvUU8fo
jPzJPCAHa2tz8jO+zzAznLGgZsGURiTehO4+wr6XcMyEMKQJHRWU47fAQje8CeyQ
s7H7F8F5Z/lriRKZ/L9BgWO2Z2BQkJl6oST5769R9uHIJRdnKeEV/AlKSw1nw34g
DXyZymIEsYdoDj/7rBr2RxWADf9ecQTTDU84Mm6qDBKP9fwCXrDCtH7ejhaJsBIK
FkxxnxeOlsPZRxOCzNYpSNemlOPqAgvVjCVmQ4vEavAlPt1ClxVZXEmtJanEf6uB
x9wA9F37p6REh49ewXf9hSnKfwzufWBMtpSuYbCErzCXYm7JgLzutCX6NE8t4PLt
8Z0qtyiJoN1+KypV0DPpm3sT3ZIh2S7OtWIBKM7x2V4y8eTA79dbrznJHpVU8KTv
eeLnV/2ppJAoa7F0vHsI3jySM8aVnsWyTBy8upWhr4SjKFi7bls9pXSLnUYfwKuB
CC9BHZUiB0xB38nH4ySM4+H4uEIhPkpLZJEEHmHf2hNuVJw9gNShbRo6VUmNaLW/
VQM1xVmL/1UfbICahlMQpVbvRq6xYvBMFf8tst9KbvNsT2CZwPRhNfW2eejF3aIg
IoRAKBJeC+BN8qX0jDp4oSJLIr8Os0M72/S7uCcieedwoV7tV5/H0BXQhlizKASf
gGLep0wtYn34Pi56weo1BCxouI3S521bAlBBNHEMddy2sm1fPr6QCgOhoIeEldTu
YisY+Ihz/wvG9GZSr5TYHeP0LzPLmo7VAKWZHqFuuROF3CKNFiqS03zPpuqAuMkA
ytsfSxxsDliqE5/f8yqK7Hsi/VdjjcE1/2+zP+7lX9Zjh9cJJagn5zx3609F1NvR
dcZiFGAIVkWKunPzBtno2ersHAISOypPi7qMa6fWlnKUsu3uq0Nepg62UCFKRj03
OTNdgDqbiibWbHE2zU5UKoafDgcYBYP4A0Q2MzdeHnkoP1qSmpTLosjSmGJJ/5x+
GyvXna0VcHCj1PetUJpxGhRSjevhkCh4rIP2JktqdZBkaey/PveEW/byZDyJN3J/
VlgW4unBlA7pRkGGNrCi70onewH8yJd93znfzQkdJ66kfzM5fHTMH8jeL+yWkBV9
QeksoCgT2gVXXB+TOrL970d7DM5OQ1tmOR+R5wLChLVeOOhi52xN0RA92hfjcJYl
S69555Df2rI4uMfF31xSSUf6vzT5hS7ob9vH2wGCvL4dGRARWHR4Whgk5Q+CDfo1
1EU5TtzoOLYO2gZ5OhRhzG8qUQfpb/nfYQDwNm/QVd8aL3a3436Q0+MvUiKVcTyH
TKVbA6pg8E2NTJv+pz0xLvBys5i2IgfSZ0aHG6R+CrhaRhoaD3LBqs6y19nhGKF3
uYutNBqkemBDx6XTE7UijFgqxmQagLyrwq0wrYTq/iDyhM5Ckz5dJBYxah+rxqJC
hPe7jBgoxHGFtk2+rI8MFPE15LPDBwuM3q0e6UmAbvgCngjEn33p24DIM2fNAtpn
nohdxWE9ECMgUrJyqXy0h887ZdtkMmyQYCiR9uMBlDV5I2h9hU3ovyBSSaF144Ci
FABtONLq87tB6yGm6LantomjlUQIecXN7sJl16zCeGnWK20/Po5wbdRePa1S3Mqz
aeo2kcYfv+YyuTi2J2+ldjZUKG5knMFdw26b7ZoGjYXYLZH8IMB2GAGFdJn74pTP
ZPZsE0yJ5NZcT+N2mbvOiYG3rStESwtJtxWGWyj3Pskj7szpcUt0nOz5Gpa/uyFj
GzM89nj0ruy37XvGKGj5on9CP2SrrcqD84doVd6I3P45H1UXFAUtJV9UlkQAyjbh
j9zq4AiUGxn5nGhEP6IfjP2xyLMwLTjqIpZ9EVRtCUUr7soBU8M1Xi/cqamP/Ct9
zCsFJmSByQvmThyV0nKdeEKg9/DUz4EkJVAOkyEa91QQIiNc0yUhBSC4VUHqFwOI
QhOHLVOLhwMkLb+xeuBwJ2Zk6jl8AMahYIl/tHHr8kAxZp9CHPNMt6avtIjpr9hS
XQ8tKRenzfFYqz9TqmalmgQ4kWtesV972O2L5KyBUTUXlYqgkl3HEod+IbpMFmIq
sm37/GfmujzehPWg11qdtT7OlS0BrXSXfFKIWXQmWC71u80Z5O96rjnV5SO5+cZe
XnxttZT+XlIDeQRTsYXszYQbj5yl/PRz6mC2gS+53zgZHJTN/vOerYWeOMVqkbDE
8l+tUZuQnvUIO9hOMy4GyPzUmsoVkMPGsSRg/70AuhRaQ4/vy2al/lIqYxXjWUTQ
NBQJ5cDOrGknWmc4iHVSWFfY/uhSuOLvfYH2foqfmq4fEQGBZUiwWfaznU+9k6LD
Yiic97oIXYZBnYm86Xt3Ip8BvP/HtZoj7ivMD1NUXXh1Xym20DL6+Lxdud5LhgNV
kOmKOP2IxzNSZPd+LL/4rN4ueNkaNrlGCduFznxEza21I+4ZVdsQVwC7750/cR5Z
yvSMn6/rKYCwJKLTu9iTCbsE9/7Xq03gUerkiRkrsQOJX9Cn8HbjITe9j1oLk9Ik
ETNLFZ47xwNvCoJHzZdnIkXR5U1flRYvnOKrljbV1jA6kMBsal2nNiAcy2o6+quA
SXohhOVZ457qojv7KmKX3ARkVNAxHfocC2cVtGtOl1Cyx15quOYQ2sLZ7ZT3rqYz
F/2vZU+zdV/DNnb6LL79CZXw3KWbcupUD7OGoK2x1ePyM7jqLoM/Vxu3BxvAxqmm
xwRPHBw68HV4epVRYLg9js3gcdV31fiIYxznY/NJpRcjpwwgg6mBGBsxf5La8m5Z
ZseLPk/S2XwArrS7u43Rvv47k2lzaJCSbYdop2nvfRby8egY06CdXBisAoRGdOf+
VbcDLovbIVdKmmIDv9cDln+LpvpxUcgbSuoEd70CrKL9rUACen8svDKIEz5sgUam
9FROytG00z4YYj6YSdX4NKAkO2K1ffbvfovkEGNNrd8tLKqEO4RrONRX1W99JJl4
C/ccxWq+hbFB9BOokI6F+U4PWn8b9142CmxUAzeTVbSQrmur8seqUghzUbskuh/4
kqznzAnK7XbqWiyiNDcZfao4fGOAQf4GTeGCgKBT91w1D9AVC8la5tI0AnFBT0bw
pIYoHnTGGW40lPoAolcRDKmK8XImkDRkIJrzqITPIo8TEvt3IY+gDtJ+Me025JDS
oEARksyHL6kwOaXDhghDRXUhLcuxJXOnsYxBsE3dUSVnNsOO1Jwt9FxbbbA/9SKe
MnmAgUos3Yj0YzYFu1An/m1Xg+B+KowMDDLCo0nv7sJ+S08Yzcg7Xf0vRw7K2B/P
7TfnVwdyeLX1xgxXMoAHmvFIxS8N2woW4ouoQb8NOTdo4elmUVLiozgsB/kUoxCC
PhF4Sh32lKRhGnFaR85z39HrWPUkE9v8hjV8N7YPYj7Mg3QuFxw7YqtApSVvIY8B
JDiUDtWIjbLQyXZfWiOSV2+KQcHslz+huBpdZEyWqMuW7TRmNo5YVz9zUzGefIzx
+HUZo/o95FRb8tLeicGueX+l7OMuqCuZXJMWrJPUsv9uie7R4ySy3KTcwmqvs2DB
/6vO/atsPlxuSoENrAFREpE7uU8AsIf4Rjru3VNkkxNjzZ8fajNBNNOLYIv9K9Fr
zU59keOKuuDcOeBZkXD8tT38rscCfElymwfj84UyqxDx9Dsqi5jjsCKi6/mvKQEG
6+YVdM71/jmBVbliE2SpnGdOdWfC15GzTWV493ZaWTkJVscBp0YW8vW2iy2jP1xJ
EixZtBI6FzPyLbit9ZJyuplrRxpDGkSDxPaJLeEZb6e08sDf3siK0JvxKmllDCy8
UH6cFplxOCQsOwqtcQM1g7Ydm8pUP6Z+TT7aINQxhi7dFrZu3FOqr+arc86F713j
9feSmFmw9xcQS2PIMfciriU2jx6LYUrUh0Ac5GmBNblOT/2zNPxS+bhdd40pPRKE
SFcGp9GDBG3tzlEsnHGvIjJ7w402LcXvucRFo/ga//5aGxy3R23ZEm1/k0/S8y/G
wuhcyhPFuRcjFPDVLsRpMCxCHIznOjhe8vVpdooFMBgs3g4Hhyn4gH4ohBaHcLNP
ZPba46+egflCjMEKp1a0Fav1YsAZLQt20SMYO4ANUFxRM+4rt8sdRb4Ujaly72Jn
UIeWynAYKJZyPPaW+brCgekRBLMFXrMB8Ex2HYiUQ8izVvfCSHZf4lYV7jv1Cow1
4MCOTZ0QWQ2Wrk9kQcFF8otE1ZyqEv2qwpp6w0VMm04ikaCzhnXgaA2frljoF7i3
/8XaBO/jcnQ73vDjX6njDCfJEsaMgFur03OGfKXGHr52ob3uhRm46Nf+IQRoq4F5
j2ugf15QLfTlO+5UJRHSYDsADAbx3EqYj4xguWeaTbysveEaejYaC9TaJDCKPjOX
uiDtnl4mmZour54vtEIlRqQZg269fwnlctfS7p9JrXLbVXVahyk+Wcz/ECReos/Q
6lsQwfzywIFVgIrk63JcJYLua3xUjwzeFGhJv1ONmLFUbFzHJxtfD/IL+Ljm0Fwi
Ia/LRblAxQ8muiBVnC9rs8TQMKPGWhaT/rcLbTH7JnRUpU9EhzuVX8ZxUwrDgy2t
yhuT+qnzIqXc9YSuozGYDzT+m0DVQQg2mbTv2P2Mhu0M+99GHyMMM3vdZtpJqDDf
LkVxi/2ioSi/ma3va7hY8BmD863jKsJJQ4cr922+vDSg+EdELvsVu5TTAIUPBSL/
lHTZdv98Rc4tm3YFnC305x+uWSqBQ5Kntcoel/NlbNV8JO6WmpR2/UFhwkVrUIJA
+H7SvJY6VkElnadva7+kOfb7s+jSj9TWH9ErtSgvZG7X2wiT1ITilddlVKUaqGih
VNBvG9La/zWb75qyZ+c8YLXkySyavqYG0NIdzznEeuaeTWYU5ibyG0CR9HB4Ul8j
0V0K0o7rWGqkvkzHMqK36YPOZTKL0VJEONhCmT+5BsJZD8AV0ntNUdOR1BW03UfV
UhAdpJML6BTrseuDr57p+eRZ2eKIufLnFj2AjFIgqOmd5k9Vvq0vQYxOiNbyzKX1
ErB4deNjdaIm5N8m9HmHE8N42UtH8uT18LbREdOumd7hpsTzbV2/QCbQMVs50kgt
oqhZDSuR2DN/jcDmVCeaCvcKGz+Z2nTtjixI1YlVKu6kKNVAcMhzD9dXZ69ga1rv
tiTK0xFcAGtEKXzcQmBuzwwfY42yRrskPaQ/T48eGWBSioNVO0mLXeQx7X/0iwgU
3b+leS7W13UMYNLU+37ruNlUHOY+XvUdRQKcPHz9ANEn4x7cgAmxxcYRd62cP7pp
5aldseIJw7Tb5WJyVOfCz936RSVb5Aze+Djzs6MvZMQCy7y6YIGzv8JikijLnJI6
tSEAQZz8ZMXxyAB51npMlfHDLcZsM0cwo6Hs2r9vpseIA4bjnyRDkXc2w+OmF6Ek
BRliJUW3eL/mO/6ajY7tawTZTCN3O3p0vMMM/WHcb7RhiIEllJADWyu88Ll9PK5W
iUBs1KPDBB3+ZZkLI6I4GD9lAf2QZmrMFLnLy2mocMS37acBTsPNNBo100Bzf+YC
lJo3NKVw/wpE9b1y4AGLzbn5a4yW6Nu1xGteFDVSrLUEVMGhksmpq9Cd1d1Fx2tE
uAHxBS6juUL7Njw9Aox6V3L+GPWrAxmokrA5neu3TvgbcazSRmt8yh9zQxvRoaTO
d8FuAI6GRhPIZHJop9P4hBUSOLVeUPhknay3A5M70NA213HdHx4ZAQV7nemgFE49
kZQ8Huy2lXzwu2ypCD7Uq8wL931daLfu8VCBueFy1lTZvwgIATl0DNQu4JOvy64W
1d2HR4Krg2r2Mi8dVHDo3NyfbT2ImKPCySWLOMsJdG5DcJAbWJXnDVJ9GldS93xp
Og6kqFGkrucstoZ8fSHw3shgxH1n1Zwa5oR22U6xVuhaqDcc2yXt0IKIpzwCwa1q
M9JKzGa/NL9wJA1OVnjARASjsj08jj1rbxUhRClFVek7eEumQgG8isnlMLQuMjCs
/3rwbtSLrxZQGXL94GUJbtqUy6BSCpIPixapAMWvCXeLml2TqC5XEOhjqnMoFuCz
ETf/yJCtld+pTUXsPGl1lYyWJw+ctfX7GfkO5Wi9zJT+VX9lldn5dG5VphzpggDv
HvhZrsi1M4LUxYJkWpcKjntKgTqN10bU8IvB3CAwbNEjtiZvzt08UppHRs7vV9lE
FoWqGQhOviXKznzUSGcBrYPC2BIUNUx+Sy+QdHFEimgmFM43ajRJlqhvkgQ4+iXB
MznaRo+Kx78grQzgtMPdTXFxeuKp9G8qBsRxmWoqpvCJE4qCs7CybwhH8OzbOrBr
FWD8z0iIuvxA6OeHdq7nCTr6LCpIHr3xCAVJHLDVML55/MEm39/CJVgcHZnUcrSQ
bsKRZAtxyDq7aNACkMfXAVdMohdLLFPXb/s8WsJ0QJoxLPbK5bTaBnXJ/o9cxhVx
Z1018W+Kamv1UgMOCvAFBy84nyhHxGBbA14Jkm4dtn6h0M3jiC8QmOO/KlJ7VC5i
kGysnrEjegYnUhljB+4RX/fYBvb6tteF1duTXBsILpkh8gkluxsyVfP1/6I9afF6
lbc2HT4uZOezfjnJsDTBZwlkNFWMnOx/NUqu+Xs2jxhh2+LRueezVlHwHPEKxUj+
sHbREny6tMh7t1MCgjLlq9ctMc+IIgVi4Lveqh8rM4hZm45bYzgGL4YW7B8QOM1f
hBRmKQWCoP+IVxZ7H43wwTNpWQUw0vFHUaBy0Clv9Nzbg3FzcZXiTVPkVALazhV4
3WeAywOHzjrpR47pY5oCPr4JzTcRYLBKU6u3+uFwJWVZ1PI0T4So1d70a+1YLa8M
uZlOrOeBKoG4VkltiQnxseRVjMXHXv5W7BYlg5wtv8hoM6hnYWvtkQk3N8te2bcr
FfIpithlJ8h5/wFYOgp+DNw5EomeIHbgjzEt60pM3fPVdnNN3hzpo9YJTUrrlsXb
YREJn58ur8nSA+UHlFV4bH+EWDPh6ob9ekb855uJSI2DFw73DKgU0fh9w+KixJ/u
UGeLzNlErITm4U5lCo7QwozjjtuJQZSh4TSybKTkCJtLDiQfm0xAsvHeCtaZClQB
O1Jkl8IOshWd4jqH6APnrzIzy5vJpQMOG3Y0bXiREPP1hg5exZibxQ6ghiyyxZIB
NELEKrx+iPqpMC72UkR3k6Y2Livp2ZxkEJvz3jkMUIN0gQma6nce5zEzdtMty62V
fJCfYvLFOVpdTjCyIJBWBk78tyMNEWVtSF5Ad1gMET5IjiTA37Y6Rwl3+qyZ4NqP
stvmOOuJlGHiGM7I97EMwUAaVFNyqomuF/PDpeNp2C1MK4N/8irydDfFiYRPH4pK
7rQgr4eNOT6CaUNo58QzSle5UsOfI4ElpxzUlMBJnlZp+i3WsCyoqLr2vnZaXlOs
Wd3Az8asbJYI43IO6kCyPikejkzHnG7YuuoFhrYQkVgqtC5WiESvOu6nEU/hz+TC
H75G0qL8rNsr8tGTfeOXueF39TAwKiYaqJzjzX6iQKb78A6/RHjFQMQRuYx/XWol
yvVeBQ3Qxcu+XCVX2f7D9kaHJ1BlQ0TGvyyw4Z1YeCJc0StNctr5BEjqn9rxvxLd
TdgDi9zQ9/NY+9f5IftIkN2gby9DWqNQybLnef9FxrEWXi1fhjNs1JDzmkm4RuLc
wb1mv1zLrWZ4v2lydNUNFobALJy81tQgdBeCEX8HlLlEXdrpSomM40DFmenvS9Mz
c7vPootxwXJZ1CSezcguB8OTXPBW6EAeNk+MaC+jjFWDh4F7QaE/zgU4gLr/MbLS
cj453dph062CtzfUoJePZBCoaqaT3t+aeISJDCgFtTkkqdkt+OmwM301fhaCuzLH
aBMWPep04i00g+qym573EMsBgMEHMSDKqSIHHIeLuIMUpXf328svp6Gd9cmQMXpL
jLcgp213QJT0aji5UaWD7IwIZA5yK8klIO2sMtKQ0NDmngAiumrf+PzWFiULJ0Wc
67ckq2impaJ4JK0WUrt8aSzo6A/6AsyKco5JHiZFcC4RDbkh17GN3qSUaCoUt6m8
vo2VP0rfQUy2FEVi1MYBRT5pJFKb4vubgfrryXDaKMnazjU6KG8tjU3+yjcZERKr
EJU6NBnsvfnOx8Qg4aTLgChSWG/QJtH6qq9HOQT+oDhycjQo3OkANXayOinRfulX
2prlsQLDHY+HP38c/l16h6LDKq4/woN09tgH+e5G+lxacUSqABWonDRda2lSLOSv
bFtcZX50bGTpSQ93vQUesdt2BlRJ+n5ngw+XQBny1LAnvQkHUdJzMN4jLA5EXsgT
0a0DZZKzPJwG3L1uJU9TTsqDV2pxjpraiOANbAjwd8KGFNNekutoXxZb+JVyeVPT
xoUEJg+VuQEUxtJQR6vWNHPvq1MnmiNO1Pxx/UcK0Q2ZE4NSEA3hKeMe7yS0Lrld
9fCpYrBbu11yUoCbh4woGSTMDvNnxKrOhrxDrR+t7SBrzun5itnXCgFq8z2MxI99
fmLcc1SV1aW4B+59DqATu1iESVKvGdEAAccQHQ9TzAkmv2BzWnM6Rf4WS0v+zyR2
NCoO6eUtsDzP4lNp5zmAJ/q9qC0zxksq0+AZMnFmxnvqKFWHPs3+TIEfD9DAN5ED
m7i2lOVmwOjtZvIzuUjB07wyg/eAfHASIWgRT/xKU+1cBQ6/7oHzlIReCCzvMnPx
Gt9SDdR6A3pIWsh8HmZ37Mado4u0QlPP4HeakaHgsGKKlCVgCMv/rWkX+GQIEG+J
CPhHy0NZQwGh+rUWs79w2Yt5QPqyhrw2c8bNOrGlUp7O5hE5//L26Hn27hFuDOdh
kDvvYVd/Pybw+NkHl5oYuihEtveEqPzBR441Irg/ZsPbJGGXOFPh8mVfrsMLYnZ7
M9BdnHvV3ZRz7IN1Vn+7WuTs+QqFAVUMI4GPCRnqsO5xVE3jTg6tZHgRFzK4ig2Y
+0hzASBQ2/Mpv3bZ+1fmvVPohfGtMgjjORNmDvHE08pxDdudWAj0+4Xl0KyIFO51
gQkahyxNctp3ZZ0oLBVH/HN2eQmkpTlXOeDkQVerKYNzTvZ/bEOhpKqKc6MNl0Kx
kkBg7heHWT9/wxElAk6vDyqsND/REf/Qx3rtbZpOhI4JsB8gZbhhenOt7e3eTxHP
E4gvJ84YJiuZl7XgBA/E93dU2JrGY7MMgHq90jqWsYh7UnEIUBXFmPwx6bvE832l
Pk0WjAHbglRzzwUc3RSu0W+j1Roqzhk7h89TDfFbUZjuG7VsQdNvxub7eefACT49
6P3x0N4PlQwBf2FWR8WEVLAVH2DJT8KAdJ5fP4432HsNTQuZHoha22/AJzs2c9/D
VvPbH0zv3+Yr+Luvd4bG6PSZWCS+wwbfYYA4ZEX4KZbCELrLCGAa7W3tWJKXFQZm
AHuYNuOo0ZS38wCmR6hqO5sodhho9evQnl1Zy4XM2Xcz4/UPSK231uzcWwwICDbZ
H5nMhlR92TlJHEXJ1wcwqML6sjmh7oyeaR+uOxSM9QV7PyZSFfJiajisEcZb/ukq
x9TruWtTh8ci7Nonj6pxHQEol90Qspp3gComUxgj80El65x/JWPxMsqri6j1XQjE
V2VSshlwFosDdS5osCe5EFx3m1rFbdpp1KTjhlNPbR2U5H9aHf1rC7Hv/D4zTMxB
efLW+y3oAx1wuzk5X7lpKNQtOlZp+UKuXnZoKfguwXhYhmA1uGNQ1HVC07qEj0Tc
LkaZ4qc+X490uYZYk3ihrlS8e3/4flw1zo7x0RQcRHVsjP48gsAY4mHikJ2NANTA
RZ+RnR8uBK2c1W976jO4drCj7T2djkz3XfGDvKuYVquzcxjtuBelNqQycVE+tgTK
Z8sVSLJnJHB1LL5zbf189DHQTxuNY2i9HTc4GAIsmmhNZIznm1pOTINoFkIQG4yI
SKObvzGI4+EP4dG+M6v93ApVl65DTzr55S4+CJ58lXbJvjIDSs21un+oU76OLPqX
f7DMFL7nmSsZT9U9yTazlxnrsTjy5dncokNkLTllFtGdpZmHEPeEOx+N+gV18arx
6AsCgH8RPFsfMQv5LwmU2hSTI9y7qYGc0B0NeWn73Ki79fdirYfSptRRgajhdEay
KsF0SNZ85Ci6aQJJCKeV9/NCtKQ//cHrD4Ctayi2NoUYqEy4YVTaQCatpuqVa0NE
kIq2sPczJY04++64zvLNC6TruEzP23S8FsrApWcxmpUEsARyhquZ3kxs98R5jkzX
p+Td87zdrY9FaczImK0+qngPW54JcVZRQzOoY5tIgcixypBaydP/xqA+t56x3xwp
fwNbbsjLZsk+WM737sYzKOLKMS2xyxUY+y9qQtS6XG34Pd1tr6ZFZ5n8udvCjbRJ
sb5Pv2y1dSu3PBCxQvDLgNvDQneaXZbkX4MkuAUssHzU3TTjq/WoNR7LmlKAT5di
319BTadLEWHfjq82uMqJMJsbD3VaBIGvrrE2tINCPnSADGi74CG3bW/tKh8TQzMb
nN6I/iQ6ibfYatXtmMz1Oo9DveG7vT6t4hiClyL+wtgqeFMVtpmQBKAZXojCPU6D
KMmKNHQIqdPNqD8vR7U5kczT8PN8P8WuJ5FUXqR3CS8/+XrmjYl68hZ4v5a3IFYo
03SfJGr4QFmF0kCr3KJZcqqpNeKUcB6O6d2tAH+VweJRQuG5DgzPTIsifrQgO/8y
dxnjwF6Mfm34I3NcflzxauKf0+MNYP9u5o6j0wGAkN7TU6hmv9McULg5gNL2QTum
kIPgZW1pQwYWLRIv2T+NR2wOeJbF58ckz8QgQllL1ANfwj30BFARq7FBeAno/oxb
bM+3g9M0ZpgCTFQaulSH7QWpUnz2GnYRpp3BXEZ7j6iMhBArfg9Pumsvu0jvcXgG
namyvAD8gImFNoDMBHVOURsGPHT3ymkjb7I+KawbeuMDOGPJoRz9A0+L2FjW27YX
cx7DfxdQHK7DLHMGWOQD5sPTjAECJo7cfDG+dbQ6SIIvhePFLH8+4urXJRCz3Nmy
FHbGR7b6XCJcsXal2UrrQ0sXs+ThzR2xNuZEfh6DqMAY04cL8ObgvW70HjV4hdK4
+i/oMHcaFJUEIcBwqAGljHqos3OIC5fzjrLMJRohRQsT7MPzHuyqh9uB4ZeLjHLY
UKDhs0GRXiwtRxYp+qm+zWztnMhqS+qKbwTv1fhzaaux70CS8g5Pyn5KhGy3lhR+
OSUXzfwt8/auEac343hGxi4bQ38mLlodG1kCFtR5w4YTl5iivJltrBewq9Izfz+w
yCzN6xJ5oNlWvBTS/xFcl3DAAmqRs2pbZMRFHpPrbby1edVQNDZSHtkhi4MroUQ4
0ABzL2Z3ptRCGoBfqj9fF1O+cINFTPv0qS8NGRh0k8//qRIWYao3orR6rKq03WiY
akThJwEZ7RayFfHFWoqYRiGxBLOBpnM31gNwJ5bQ2Txs208wEDUMRThvLhioRgj4
E3WGIEkuO2ycARLzk6mpaLAt7GH7iNjfqeEvudNKlbg+6zUn/7zX3NxJyrYioiPe
TKNCLrCtBGQuDWkcAijJJNCqKIJS21ISNp14X7PTpKQxCF9tq2a9jgV4M0HfRrMo
pBz6ZBDVaF2aGYLTiG4XeoJdC9rtX+QeObf+p6bZiHbNJDeowh4Bd90Hppq7nMz+
7MBULqRjJjMmukXBgjtY6jId2PBemSsmPmLhwbrb4TTt52AaQ3QSd0Ft1YJ2p4A8
Qa1EUof3gyfuaqZw4wXn5bupUO+VFb10d9fAak6XePYqNCYQ5tAA73p/FwVDbklM
arcLBkv4vGE8ZQJH5X5FaDZ+950dDAa9BP9uqy6a+Pj5dK/8dcR/ZyQeJ03FHI3U
qpgBLESlP8GFY53hhd8b0hgU+3glVl5YHeSffwCdlCH2ubOnBFKveMKvgCO7poK/
7IE5YSVYjbsPswPgrA3yj2vAZmiuA3ok5iCghG53aVeP/UOpbOrmgBjdylT9iKi+
RvwKqsNta40aQPdsLlRx3s5/IwljS2iOc7UA+0XeF9TNOov9ysqpqPKd5NpOD1ZQ
ETIDIRL4g3AOPS2aLoCqy/2JHmyN5zIZo0S5aSt8bF4bHeg+QDCxe1t2le6pwzB1
HhspXEz+vD7SvJoTiI9ZCk3YcUh5/K//loq68Ex4HGYkm09NilqjXh4LZvKxru3S
Ir67xwyQxsn4FryjcAGiKhFUpsDGP2MKJT0OKhV9RWtd3KKUh0IUraszPLi3qeD5
lz/La1/wGdrotUzMJ9mD5ZjR71V+ztxNyGPgbvW2BfN7h5zF7KBawQFgbPTGvDVE
kGXxeGTSdpaRDVyk1/dPpo2uBNJfeOzmSSBRJZBOJGSFFPo2ey/xOzEcIxN5CcGL
qQtbi/1/PoqwtUMSlWbNBxANuOANe6AgvDiJrApj3qs5uzYBEfTyS290CRUYoCwd
t639UbW/emSpy96oY0c7h5YumY0icvIQfbBTICz9fXwBrz2pnj4xG+Ua5R5IOveV
Zsvd7PkupzGTgCbVea3RG/YEff9Wi71YSRHaS/LaVYX1HESKYEBYmKsZvBc6y2lo
qkd8g1fpoZ3f5zZaivAMgNDmdaSvX9H76y9g5CbglsRgQCK6ja615kfOJZQDRwCM
ewt9lID2L2dxyFGbu6uMVDoSECu67vtl/oVuhhLu5Z3i1wU1XuAUoLea3+BEvXQ3
W/EehxI9MhZ49n0Q9WwaNzATUtukzuMuX2FXnTPtwtWh7TIG1RzWdt8o4Bi6Iss4
WehP0dqVebmlV7EEzzcf+Tx2UMVanZVa0uPlpJV+9RA+wSR8vsH1fvy1AovOdCqE
IKVsK8dFtMM/YgPrFosbC0UHS9k3RKDQgy6gvKMEvGDQ06RfmajKoCUip9Asaxzo
Ilyy5rkh+MAYhT6qW0qyBWSLVImuei/jLNBqAsg43x81SIGDQxSGaf2JzLfjEYHI
KNtbytFM4YnyBgxtOKwtYzjBnXmkaej26JbDVJGL1AqknxbR73eZYGCkPDNgi2ju
jLIkPx08kXzj2339tCbPZyFJ/RfUAIXCbyHeTmgdhTOzXbx8G9vNl+fXII2h+ZKU
RsSr7mw1uf2QO8K/9iHJliIBLJCkUcUFBVnBOoVIfg/czFjuW+7oDbD+xik9H2CW
x3WAmyIkhe4nEA6kUcRrTGq6jWCxjaUaVmQC5cmZYgqSuMi1Lj0kpwYZD8cAKEQv
RW7P5WuIz93n8SfPwwPnmEFyWseBdfAGJUaTI+UJO3jwS+lC1WwF34IetqG1aUtj
wTaw4mHQ9Fj4pQgRpeAvdrv+Axr+bw0nF3juz4NPd8XXoH3UKXNINgyw5P74ft3C
tZR1eyTKx1BqT+Hh55FaCg/2iuvP/ocVryWEsCWZEdRg2eP3rRqlZMrvGUi+oH9z
HJr/XNPYXIDcku4kKiW37S7OwQhwoKRHpNHybBsIF4+IsjNEMzMeAPr6swaGawA8
TTzvK7ZpUv1cnx3lVUeMixj5LQ8TQ/Nkbae+jYPG+BhE9t5ONz+o7cV7hA/3pvns
07pZKjynkoi1wkRJZU1/CJbUu8rX6lGdGbeivAVduniF7aISrohni7sq2oOFn8vo
WK0Rax0FEQMtXAUsQtCcjYvKF3e2KxyzBFtOC3AtFd1G+2XWQFDQXkM3f7EkyECE
c6OMjE67azjdoxM/nBnHnQuFCVa4u9+eakHEdhr/hcgYNtL4ikFhY/bNaWfbFdhy
oBMbsYuhEi/Qu1s2TmcXUt81/aRJ0HIdIKaZUCjb3ux406VwmsGJEvmt+8g9ZkQy
ESpCglmJt/QqGJ88sjz9D3LXSniWQKKcCjhHYkcvkELO8nSAt1UxnI4ttCvG/vUN
BcrZdMUpBdv+BS9h0xttbya1ATamj1AY5vfYPx2X0lp37L36D/tgOImVaURcUCJH
qAr3cSbIEu5aln90VVbiEMC6c8ih4TTpNRqPjRS6q+mjgXRx4sJPRYRjZMHuV5W/
jsvUMb/mKUeqNuZCIOsfn7eJeH+2QL2f1WRE3mLDuguDMueIaVT3ridxA1Vb3J6U
MduL+SrFPRT+YBL1/lCDplxthto7k3e3Jsgy9tL8zw+RKSYaZAZD4nxl2Km75Wdf
M0Q4mUXeambZ9G3lEBBP0jAq8FPsZkIS3I3k5Pts/kn9wzvgyWMfVeyAoLNxSBs/
5FBbCUg0putr709wt7tWMQk66RDcx+gjjVBWyrS1PUUJU4+OsA7mJIogBD9CiKu+
V6IVj4K55J1OR9d+zWwGjG/9aIuOS90dy5sViLvIhgaTj+mzBOaEqgJpZaXh4RG4
4u5OkCtxxEKgW4n/btEYqkNG6T7ETkADd0iI1Bog7XfL9GmJ/5uGYs9OyyjrvNUs
IC4GANFpHJ2wlWj7Q5AJXYAJ/XaOvEjsBlF20VwBLTaZtGzJNvuQqh0qnB5iM1AK
P3PTX8Dfvc9cCCyBEupRkScs9DZWIANxfP9Z/1mVBpkFAUOSUzV0iZ5cAJmlvh4M
aHsP04cSo2nEVSy7/Do9D5TF4slKrz6aXU1DrHz0PW5Mk2eO4fJ0EfbgWdWdRYZh
LcLnsWwFRvP/Te63FcmYrs/h6BuUMEB6OQWNSAEJYGzpY16UFfmlFEsejlidGY5d
QbqP8POFnYWxjAkOG77pRHpnTixN0IVa4sSEOrwNH6ecoBssko8TdzcK58ehgy94
i2baLol7yip5jYFGksKCdGoiFuY2dqjb0QXJDXaZeBJaIdiUrM4bcJ2UBO4N/QBT
0qBWZINQplQW96hG+TGML3Ts72ONOlsDM6EqifO8cRIvo+I3C2npjE6UP92TUcw7
SO8PKlihDCwCZehnlExqPq7AdBf1ub+MZ6/o+jHInPiYNQIxH8u4XbGkhc890sCM
F3NJzOTgpcLfdcvjrpq+ogb2phge7TKKAgrifwbWOyMx9uKiG6tY65XdT9A61cys
Uu09yCQcKVwK4uyvtyze3E1xW/In1ZURGDSvMaTCu9qBctBEtSbLZBwaBdSEVhED
9XfXpmbZPagzW5XR3/n/rrVUQbHwEicChbY68XCGp1YigReNU3qHBvXoR3Fpm54q
z1eZw/oN4SR6zTqY7eDU3KkZ96bL1NAO9m6BfNgjU+wLlYxTm9nYHYOP/FsPgbhf
y9ik76rrKdzsNTIfACPgO3VOXPRbLfj5QWrZGViSnN6sXjvNDsqblj0p/+M5RSkZ
YQmBtYcWVMmFXbFQaXk+qgsv+8fMUGSONdAu1ycpiIguSbc3pCWavX0+gG+k9KoX
5HrPQzTLWWUT7832bmgfPMsUSd0+rhJ6DOqSxmDDYBFddmKb945Wub5cLjJH1Bq9
vU5xX3cH5AI4WQusA7r70NEKIn1dSrLqVqf96x8iiQxGzle7E+dowWl+J/21iV3F
J0SsPqqjEHzr4vOFtPG0HOma02kxWAy4zqX/inqLRf8sYKG01xAyQ+A5YhqSTTZa
vlyqAE1bs+5uXLVUh/8lvSQ31q/IuARHGEjJsopcFRfpG2L5lXke8ka9y48wSWlN
UYV3zRNgunVk4RsYIrgaYPzn1g1U7RvfLOZgv5QyKfGtXr3LjCREPakR+AIOd9vQ
VF2/9ljEg+W6EY7413ezI4TTDk6MyNrmydwi6CfJ992T/gw0IwXUR/B6R/xRiZdX
c6dFHaq62ZgCq9r2lfEAJ4A4einNUUs2YkUjOCfkWj8gKwvgkHMGeQ0eelQkH0RH
oHJPhnaHDZ9C6Ra8QbR/NtLnWD2sHsPWmHZcngQGz5SmBDrzI6Cy0M/wEmkzqW/Q
NJaD+Fq0z1b4ar7vos8YwrOAnTCAa1l07uKLmaPeOVrdLHRphd+m+3eW5hvGRmdS
P7vECcLzrCq2b68wYppC+oeNQW7YYkDMKvgT5JPRMzgrsqiAQD8pnJe1swB2I9Us
Yrhst3Nx3M3xcXGxLOftFkNCNZQRMNsax0RS3o7t6coQXkepgSgYsMRlFPRAj2Yy
TMz5BxqEFFMevEzLHrEr86nUmTNT8iZIivP5OpfEG9WPOBIOLd5RAYUvWx5Hq2Rd
MVjUvPejj7llYq2Um1t9wFg6gr8VSqF/yGnSIJjCiQSEHIIlqGIrC5VnvjzUqoxo
ngFmGGfMs02RcgIkgpR+yqoKujH8S988u3EhAJOtmVCfju42h6STv/QzIQiNM+Bn
BPwSxNUz/rji/5L05gPKyvyRz/QGSB7wqri+2ZgtHnHTwzAXVdC7KoGWLyCUth+5
AhqnlV6pKJ+ziDo5I2AIsGKTBCHH0Gidp5Y0ZKGMpyyZVmGIkFopbDPucL01P0Cz
p9BgwneWFOlRjGv/kY6cn+YVLgEwIFl0LGRnerVJswXklxzpq640R8HWuCIcqFwl
OkTW6DawewP8KxNpeQjTP9PhkT9F4O+6CTEZYF7lfuKADpJOwTM4KNz+qsmNvivF
WxXOm2E++qMF/VgvdDNSCXmlgc2gSrfSg6FFbdPGN3vlSeEF9y4AlQSECxOntIpA
lwMJT5eA7NSBoACpWutCduXO1XRkzYbAW9QVHGf2WX3bMlLqP2QtPHWiTsQ9zMm4
ypPNZyiVdyu4do/npdlBD8m69Uqk4iehClAeRjQRrmsh4bwhdl9slvqE+k/6//Qz
t/XAAMFdYs+NWSwr8BzeEORNsWNdG8CjkY7G8QeOX/2f5yNkmIKQES6eoBB+R98g
Rkq0ZAsejcQe4TWzoynPfiCQfz8qqxXywLLyQtjrNFsAry8k4txvENYbhXrgbRzn
F8C6vFCIi7pRpzW20gZYcJn7yHY9HBC7lZoN6EOOzJZ4NFvj6M5T1U8me7JBakRs
3+yj6aaBd5MQazrhn1mvtlz719dxkfJdLQL8nfe5h8HZ1IYVvwvJvyVnRt6a0Gvp
QZE57v4GUx2WVjThsDsVod/0/c+S28OebWlUT/gEmCvz560aIcrjKWTaGo5j6zFU
0dieN/cb18jLvBhRPTsA0cbxBPBiE2GaWvcADNfBW+ClgoICkTlgFM5W39IkxdgL
1zTsCDBrYkr3ZgH0FCQHSFmNH8XJpdUl6ISHJCny835QYtDGOWtxJdmuOdAzaeD6
D3BRDzuczi3wwAPvdmnEpiKmM+nCA2NHDB4r6kZUknU9rj2YRS/5s4Lk/yb9H7xo
YlsC+ZTXU3lEuHTol233bVSWrUcMjUPneGeEDeZT6Tr52x9MtY/Bh+w648gW5GJI
mKtBX4XnGPgfoz5cMCQ/ca+boDBkOsKrBk953TwTIlI/8v9wx8jAod6BvjxsOxuR
cOqZYksGiS0LFp1uD88JIceA7aPcyW9jl3HCQRSKWZdblYLbAsjnRNHD1ok6at87
gJzYAueHnqsQTKXHKLeL7R/2bqjSOcti97L2MTt8SwhslOTSKG6U3p/14n9AfZha
ZDl1pi+j03Wi+NJ22LDKrnzUQBypa58LN6jVP9tfgHgKumoBy7RXQwrQ/EVUZ/aH
TeqY4S5CX6U0b1aOYxSzgh7zd8tHnGNua0e7PsVBc+DAL4AkFvyrqRwP4pTsm4Up
8yhaLavbMgFCRciSd6e3EY1zJiZTN5twzVuLxKwhy0YlKk8ofh/RCPhAkNTuWcaw
wWTZQvMl5CMqf5ObapNzUSq9LOx+kNzw+aulSB8JEwHWicyEwtrv/2o/qeUpehd8
l9+km/pQ2en6uS5o3Wm8xWeMKSSatNjugNLNsqtLDZaLohZxILosXPIoemKWJ3q0
GPbVoJkx6/V1L80V8O5UmYYLzZTtECsDfphovgm9DCY2DP6mvbMp4FE072TPIg2M
YizRnge9RHfR0l95HjGMW1M9C+EQPTpAw1vF1piNthnANw/rg4qqp2WWFNeiua16
ZVyy4qOE+4HO0wn960cS/kE64tn8ImgSg0pMYYoQoD5dO9qIuxlpwayYo3Kt7vu6
uO3YrGB6Bt3rJCXlfQeS+8JU2LNg8xUa1oLbLW7mfxOU/NPP0Oz71QZ8QYNbYy8f
TOXh9cUg7YkX90lrH5OvICtR5Oc2lV9gW8v9AgTvOBFh2pa48wtIKTj/JuqwTEZh
0iNWzAzmRq/Es+UNF05y2RTSM8gthvEfh004liGvyIPHGd5UJuq2HWe1hzsl8zMD
ejAOnCEq3Tw4Iq7VvYwlBnoNszOCeBBT0wVEuKNnP31hNt8uHbfF5myVD9p+VI9w
aZyReJcd1kIG5IFW3PvbRO7TO2WVh4etJPed+CwMADkZX6x8cFAzRtcQq9lbDZZ2
YrAw0+Wq67iEmyB4U+65V/3jkL3T27suWTviv8KDamk7jUn9SjhU/sTxX18ZJu+t
To9GaK9U2vzzI5rnxMb+G3YG4GJBe35KD7P4YRVHPIuOKm/URLi81+tQVTB4JXGd
miwnlu+Oj5OAVzxaqgFyyM1zkFPOQpHzMtQ6LQ2VaW+KcW1bgkI3+8TBb9UO7uBD
eRb6r634D2M4hcEnc6BkBcjElCS8oFnXhNjFWGSJ7JFY0yZrQ2AkSxvG9XQPsim9
2UOTeJWx37/ny0Krc1jHNhFAaa39R9ksVXkByBSup470gyVCdooVw1h1CWCL9QHi
BlQCZD1Pyf8OqgvUcBo58H51trrIg59CcdUShlx+LA7y5C+sRKTvK63nieqFL3T8
UpYhB6jfzRP97gVPzps/ITlGs5Ksl+D5f10NfVRPygGA+2WuM/yFYLJUodpsNRdu
erfJUQHF5rsAfoANzW3dkl3vxlxT3SUlDQjjepC9n1oqSFSE7uYaNx1b4NOhzD54
0dj/GP3FekSEvqFe0PGhka+EiPgwpR9PUhQy/tozyRw/bsoZ76ZjntihDaECaVRH
VaBSonnJ3BEDr8nOP3aqDAwbYlwpNyMn1fYvSCu1PqQB9EvUOreiHc3z4U7h8RIC
4v0Nz1m7p0KSBi0w6n01I17SO2ji6EV41RNMTGoM7qa9x82QQBc3cGJiohYWtID5
wcmDU0+9gnnZb4Wh+ZkHj5lFDJmPuLEE3IRz8/mX92f01Zwa7zzmEP3IVwJy0sbX
Z/X6PriBQNxehqAtuzEE/4jZk949lHhRmY1pKNSA5nkjasUOd/LnxgNG1cMG/B/R
slaPnFjQwps6UIkBacsA8ZFqNpKlZkY0iFzDPIfUpxglUmvEVq2srWJUUu7du5Z2
JhEXWftnmMQ0GCbJCrITjxJEfiV0oRU5yQXALDAR1frR6Xw3rNKVN1NFeaE5f1Vx
9MKCAInTMzrKs+I+Azlpj2fOY0HTBtgfYQUGy9amcQXcrC4fzHpINvyAFDdsK0rf
ioXye4JnNCN5lGEKXKPIIzWXAyBwU5ICfj6zuyQsbROokTjiwO85HR+tGXSRdHBc
gfegGEjShxDXo11T8Nfp2KfegvXxvoGMvA3/tW6pyhp2i0kaBq7WEe35oPhPJ89n
SNcaHub2FWDP1KJ7smW6jjJW37sVz9q7d/HXcDfNUZi7Qrfz6Cw6xD1+O8dhlVH5
JuCAKyPz/JIyvWSDaXHB6D7zxFm6cz3hFIVZWijAEW8SUqVeiCLI0PKSWJcS3GLQ
Mc+hxa0idBy5cP7TGWBENAFQpBV9nJcIOz3QVe/NEz9BzzhFsDQOFTFqVDb7zIVg
9MONFMSzs8Xu3q5JnhHiA8uwFgCFTq2a0hGSc6kHyY2OO097sxnLk7Lo9HQw7aOu
zftZDaVbCOeJELqxsBm5aiCHd3kCbuaPZQ9UZqLZFu/2TH26dY1BAj+qo6DfpAW1
lrk4UK1omQpZHxHeohdOWouTYDEiO7nSjNzHewsra2fkhZrERVUr+GQFRlNv9xk/
xARppow56/09lieCexIH0N0T5Kn3vXMl+1gTccQ0sgH7cvnOX33A2A22eBjNNaZ9
7RTkRgQRNXLLGFXE1Ms2GQifDr1P2cFl5lQoA5cuq9fBHKci6QqsuxN9vRQL7byD
lSKSRgae3VFa3yj/r7g7e0hQOPIZ5vhcb2K7kpkUHZpGKWmItYxAjiGWxo7qJMmE
nBYUpE7PGwF5VGlcSU0SBPVyBc0ZgtEodIyDN453XByGWCg/fUGp1Tt467z3eKCP
X+lVXFNUdfM4yGc0mYB4U4RL2Vz685q9EYvWAegV8a8Z0c+vaKOL1RQYwGssZZ2y
xy5Cb6OAxLFF9BUswmGhEzHp9f894AVqPRQ8u9Lz+kuiF8VVRP2BV84tZ7BLRIdp
DToSQJeEfPPDcMgFCeKAXkefJyWAAiaPAOZifJOKJUmI7Rulq4la0EtENMIL57HM
HgMCZjxuqs0rJ3GUiN3I1bmo2NaVe1Li1pWLWMPiLMnPYTLfAKfC85Ddzr+iAHaR
e6oh4FNnYZjc3EgQncTW0N0z4BVRHzORjafoAnj4OHdW1kwq5AK6IhESpJhzcxc7
dGWbGE21ZL9J5SOjTHAjX/Izfq5ZdIxWZxRA9cK7+eMqCcM39v8/4HChJdQ3bzXT
O7Q8ffP4Nwug7bYHFeuCEqJFiPGaQCOx3WuKB78BeRPMTC9VVo+xXYK2TOskN/7U
XQhIjyxcoTeWGXtWK82fKXsHXWSzGd6Lz4h9SVhKb2UUVGM6lSwf7GcWZ++1h0Ub
xofHRA20+jpmLndbfMpDCW3bUEC4FzZmU86e38lpRhnLdIrSTpwAWZm/XAUx3imI
pX774U/+//zofRJn1wrMvw7KowhqlR5koWYfIWuCOEJXcN1y45tFtW+Y/pwSgKTf
oNf+FAd4RC5er/Oh9JK1D6FgoAO7KNBrmkPU08SjiOduYV8dRibsy27Sz3/qB1lX
Ng9bsZmPXXrDlr0BSBpLIWOjLJfHriJu45MHkE/87fhjbjaLGr8+XKh67xuUsWF4
ELveEWx3huTd0+gDSuWvxzGDHpAw3AUQGBOK4NSoompTZD+AqfOMFA6Y+LOz83qg
d1ZplEyk/KbAUfhNjYOxxHUBKIqfYR3RFd42ZriuyXb4HRJsOyvP8tFIDAQcgMe/
eA18FWZjHqrchj5969gNhCGkDytwCq4n1Ef0Nc+A34y1DNEGu7BCbL2La1tXH1dw
hdwYkjg1jMmFDlHK8sLCsdHDDe0F/1Wl7nRx0YyauvuqMY9oVyUizUWWL710qiZ4
p/jekIryfxSklG009NP8M5Q/iZ51W/t+2hgQjL9wWnc2AFEpIqD4GB+JutlZJneX
A46Qftjh+hLMAruBCr7RKw71tbDIXY5QRV/pWsvNHFPQPs9bZUR9S+agxqbrP0Of
uPAxAFtrlGX4ngNZSF16XjFumNMpwdCDkhEEx0foZoaNCwbjcRZTjslNd7t7k0Lo
N0gHxLH9ho/yK1Aj6IZAPreCP4a/k4LRRSVKe2b3Fxzrzgx6wuTMKJ8HSKjvnMWA
ezIZN5+zBmta3b/atwiZp6thmGbFChfEOoT68tVHPd3JvN+9ooRWG5D8YdMgvER3
U+02ZJ9ygPpB0y/IFPMYq2lgsjoXiPUzImMZ/ofRLMHqg/VN3wfd/5POGGbrbpmt
nj8k/v7FwJO3gvZZoqMxV1xEq8Whc8ZTcWmRNmTJBHvorZ2VaCOYuVq+rDXA4o20
YLvCnBEfVU6KviclcBRZ9XwFB+g3AYpqdqOxIxLYRiMSRUMffzYc9FAgFaMbPnRL
yKYgBIPWYoBKLo1mOPVEESNkWX4WJAp9ltzBahV/g6+NWCzcTPZ1tF3m7SE2QxGD
WglZQt2a3cT0hAS22M/6BuOAtg+xl63L3ghITOL0YmMGfzdxxD8NRtCIBD6rMa38
b8FDoSKFJEu3H87MKzpSQT0mNRieIUYqt/OZBqlwWKqlZJpSjZ/g71XaNNNASox/
1VRMPXvk04McDlLgFgYCicNHVK7QqQvfllK/+O6JS3W+TtJ/KuX0JK513zH6byCB
LO2i6BImqlsYgIJJYBQaajoWeEn4h8Mx4xnF3/elLPl3rETBwxc4ZHBMRBLGkEJc
qpnFG0kRIPzm7H1u3oCNH1d+VDUEzss+fjVudejNlQ+PShrC9c/S2ZUAQQndZRIq
b9VQ+XtkYEemVD5W3jr6fBJ1HIAxaE5EfpRQg1vuX6Xb6BWlhJisBsZaKhl3iwwB
sPIpGSQSfWmolNT5H3HM8OqJ3pJ37IKIZqExiSkTL71QqFjLkVx+t3XsMmSgDufp
vLrn8escvRjGbFKqVuFC2+YRpGUF/jetRRnSl6GE8KvqIsOXxAbQJapm+eZEOTtB
uiR6M4kZf8sI4KIPrqJZZRdfqiswxDMeuvM6YF2bsd5l+WF6LCk8NElu4ATHHbag
ARH0NCH0xvU3Ega7dM4khMixS18DAjfgrrlMcREMJSXUWLN/0HKSuwn1Hds1LoGB
InBQVdY3tXkfbUhKaoJGj9pT2fIct2XaainURV5H9az0j8zQNv43sX/FN0LmK43P
Nx2hOsmHyQIhyJhtQguGbPMTSrqRcvJjpP6LbwvyUuYHcySCSRdxCXo2Ggq4EBzw
ynWUzCIGJUnT5HpLWnrtAM3KQzlEUSHjLfugz7z8sWxuO/F+83aRSg6UiRBAWEus
4JX7LFeJzWq9umHltxz8obG8wruEuWMA3e8gKYiji2L17Cu8lIE8p2d3zXHqX+QN
DDX3WWgOGM1Gx6qXb+CuCsrxMi/NZlbbew6BAOFVDgt1KzS/HjDLkkgbsusbdVcO
ONI8x/s6SUibAIN11QFOO4mFn5HeNX2yGqSpOp8XratD6IEm6VWiK6ZHjoC3ODym
5qr5pODxdvVKarhTSyqGC/97g2tfFY8Pq6gYED6GZe9iZxCV2WZzqSCVBXobJYuE
znW6vp3Je+RskTmQuGaMLyHRqP+z3TZuRWu8ayH8g62UZD0OnvsWRNEwWrzpNGAK
pNz+Vtv3mDeTPjbaN1txNZh5lda9x6D6DQJdqMgcfCCOeVlYcU4MTrliseEdlR2G
VF9piyhE4+wq0Sg/N417YjbDTYAyjGGekHrMrtxIepdTeFof6VXWtTdoYW0tYa9I
nmBfsv9rDweef9aDVgMe/mciFKFEFW6rCFV/PtS6IQOwkoOjwj8Cau3RP3vQo9Jd
RyIVS1ljoYImhU9UrBwzAZL5Fxx8hfMVvW3xi8AgmGoY+n+EPX/T9CNuJBClwqW9
r88SOqpqMGAnBWZVDZWVjaIoSadB5jWwt7cxI9OpeRsKPVZlcsH8KvQXjHm7U+mQ
xiKBg/mpZc0shX1Mo3DCDhRD+Y9eeZ/sSfqrdrOR4dTrd6AAb7TGem1Bh/tmEttS
kLvANzYT2dusbgDDVTqGvpNp/vKIY77Bu66O7g/9DsGGzkuG70TkFKIH5hG4QgZq
eQYz6c4ViOBT0qEeCeGFFF4EVtYiL7HmtXZfQ+ScUQyMnNYU1dN9Rc3as6x23pYJ
TGTbNtCuiqeqoqJ54O4VwKjHDBTLBv8Tt+zAb+5qIhJx9EKGic52xSpT38hWfkaP
2Nl3erZRnCmboxOfjiNSf/3oIE+lzXqe8Jea1Gz14k2lzSEIFGZa6M2EK/DpE4jW
WC7GWF4GPRi1xt3TXcoKuWrqwohp//TvvDm7zsiFsy18B9ru5kXCAcbKQ6qXuMGv
Jt1ZmvTBbNR8CmzGIsMod73nJaACv8EjG2yc0DXQ1kn5KtUN1dPDVSvge4qSzDLr
RexQ0vtw/FWA29gGl5LvhVif9KOnDLfRDTeEnK2bc3OHBGR54z21edzYqZyLv3em
cGTxzN2vCoSsmBQIv7eG4mQGc8QAjbmL7j0/7nMyc3OK5fXeYLaitnG6Ul0Le0EW
kE2N2kjA+DL8jJs4nXnFij0wBJEMPtiaPds7XtGi9vRxq2AfYxEEu2u3OlpUVMKc
vtA+8or4ec15hHW29enESI7sw5mV357scWwQhbPtQDqkMhKhDQLB9sVadBDxrjHw
PAdKGQKD6CizYSJ7gXSBl2FLYRbYO9okBqtahXRkPOHVzoUmjgqdPJuSngXkA6gI
2tptTkvJMn0Up7CEohi0wrvTRqdjcZS1ZUGtHw9MC7+t4PCmzN7s/JSMRzV7XqRk
q8FhWvW4ly+WqQKNCJvLznbZwxjHSxqFH/a9Bu22aqPtkBfDEKHDAJHnM74COxD/
WqCj7xb7GNEoEG2VxIe5BvpEGNyxXCstSpxheKr2U33PmJKi24YDLkpBNw0Apu4t
kUJ55aaoDt/Pb1r1TA6MZgAdhdxswE82grypRjhw0JrRZ3dTMEDgpuEFxs4aBPg1
2wYhagtB4/AMUwVGlw2XEw==
`pragma protect end_protected
