// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JMJied0v/a51yf7zK4ytnFkEw/5jPAtVRSnlX7RHLGwuEWDKaaHkvKIas1oy0Y4d
TWT8L/PCEF55rmc9vurxjRNOlPN6avHGHH9lwd1bfbERypf7tmIaWKUv8QBbzITV
JoNRDK4eb9TI3u66HlEnJAs3uWzWK0Ts3Scc8bm08Lo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33104)
jTyp2JK5vJ3LqXjJ82z5dcqLah7iqbfdERr1o1GEA5AE1hVzr/FYHWi2C79LXiQb
577zQvid9UJ3dkjwdu8dcsHaW/SCUB6t4tmfuzlGR98uaCGRj/4QXp51tDpf2IML
q0HbmUQ9wgGD3/lbU09H/sSXvbYfpYgNHtRQAVWX4SwliINaJadHBmwZVgga8f9O
E9oPU1rkmvNfBj7P7Jg3aJtNeMdXkgcV0Y2mn+LSD+efjC85LPLkqGFWaahtStOg
5T9GCIpDopJlrJe7cg3QOJ5mvKVad0Rf+7+VJn07035YtF9gdeOXfx89itcBl2IE
6+Eip2YZZclmDcr+Y5/vfrwDH4vrby19Ue/Y1O5i1KEF545roqM3l9gemphSmSdN
toqiZhIc8p2Q5/fqrATFObwNnbzBNuvPdhFcHnZ0cuX+QZiP3LADTqVOfR23UzTE
G5D0d/VW5AoR4m9qBnmxXuKu9rxXxwscnuDAPncAAJzaVnNNg1jskMb9AcmpQO1Q
XWIh6JeNvwCLjD+gljbp8E1Vktig4Kb+d/HFw9QdrOJzH0JF/tPFv+RTwsyxCZEf
0kugfXe13jak81DfnGKD0951NUFQLauKkMvxF4NViP7CTLTwpEE8A9Q/1bPYyqvk
nUCfXEdhO4K2y/QLRKW+NmtIA9Bl/adlErY30P8zekXrCVpQoGrE2+BBRH6tAqrh
5XLMoMppe8mitQYwlpB/UB5gkv8ZjRlpqsVSYR2ebdry3qTnC8DH/LHkrKaSmZm3
NPWNEQ4rRMGGKnO17j/v/X3fvGBFPKc5n96sIOXzhgT9bTDPgG6AqobOu03XWO2k
lXyngYKcveZ/PFVAr3auadh1hJiwIEi7M9Tfhm8OWpfYOo7bpANWELeCF7lTguWP
Izhjw1Fyom27vbxa+ier8rGlpkwt3szGCPH19fg7NNoaoWvvJhJfYp40umk3Hd72
DIAkVeyVCLniua7+BKIDxYz3OASO5czeRlXML/DaAzAccYS2euJGdSR79+7057sH
CO7KhGGNN8meYqzR9rfAN/Gqub2W2bD7bVNgxuHaGKn5ksLBkxpjZsBNRCvlyT6Q
aTh3XvCPSTE62MIGpCP6eOX/GK3ErjHTSk5Y7K4kHDzDWthgM+im26A5c+O8GeT7
+qfAA3oH+V1WyeGKGysNTRCp+KxrkawZ5SJjBD0lWeF+/0GTh6YRiUxyJA5409A+
erRvgEYM0A0QiWlK6RvJwqGOKDGSEHTc4L4v3N6BZP94oizd59+ugJEoI2hYFslK
R7B9+ERmbAO3eR/Jh56fpjgHm+JnXcJ3Nx5ok1QG3gmJ636sHCGQswoLHU96IY7Z
ejoBgI9BVTcwro9KSII51RI3HZSKy+CV4vRNIYjL4R45UaIuQwsaYtNQk84QRuik
tLVUwKuZs6bO8CEpUnxiIRU/oZeEuGiTsHtDq8FB2jhJ0tXKJoD0deAmCfTmhBjo
fw3SeuWBavhsH8YQnjDTKWD3F4QzSzJhoPMlL0guXMniiVvzY7d756vbFYL7hSVR
+RE2SZcTfi91bu9KL/NHtJSdJmJSf5FZ+rIruKfW/U3zM1vFlvT86fzqWSV3uh7h
WEmEgwrCfKaohggLOBfXSb/0T1P4mx9yB4wjgl2A38ch6YLT2XFXZlwUySUJSmiZ
LnexsYNwsBmEjrR33yUBY/8v3sedcCsptSpgPQrksITyMq21dkPxskP+WYeScUZE
vnXHWb0ygzpkeqDpXRZyKuWVw6LT+XD4V9LCSsX57vFpXNFunzYKY45Ug91tKEU/
HvN/Q6ULg8rMAzsBEP3wXCwV4qJnOoCaawIP1J52VeveRwH+XOSqtLxqk3piT3dV
odjrUR+g4M+0wewbUGQimshiYeri8SmZLNtgn0GKgatcui/OpBBhrxZcYy2tQS7Z
ngwhPjSAHRHeMXyrbEeaRtlruUDb7ciwcC1xofaQV1yUmtCifh7tcpI2O1fIfSrU
MHPYcqJPmrvhfOrzbBwDVrHweSGYlseBpJ9pIgQsAgPHKonv5rjJZ9QucLgQs0V0
O1MeN6oRf7qHbnVg24knLmI9xu0luQi/siOdu/997bsCRL1GTei3Vjdni1f0qiWs
HG42W5fkfsbRH7M2Z2C0yDFcuGzpGQS253cvmh78X/i5u4wc04r0l7FRUjaIRNYZ
jGaZwlOttqg49Eyzl4kTuFIAjQklb61c5ebUjSLVzFnWiWIHOMrJ5pZYJDL1e+Jk
o9SOojiycfCTAh892eWToR3iDD+d7KVQLoH6l+qA6nIpM89iNYzYtRHCD/+8qj6r
Fj4ZPjSTzvSAay9k5MDHvaQVR8Phq3Yty/+LryTWg+X3hp2AnIZKA9GqEyJqmicK
za4PFn79+1lyR0zqsxQgW9hLwf5Og5sPQBO+/NmK6x2WR+zNdf09p0+L+XUTym+S
OOT0q/IaRRlOripeyCOacuMrB84/zp3zTLqz82F3L9DHd0bwU4dfT5ZCS1S/cWe7
x7er9o/q5AckmwCr8BkxRwax1SNFI6deg4Z9+KU8nQbqldNxhhOhW0GyWgXj0KyO
pluCzgU0k5B1rU25ZcVh3RmkEiWXUrCETmhEy/J3QomnYdGNjE07QED3Xjp7eTg4
GsZnAp5rzNp0YZ5BASn/omfYKjGQy49PwZzNtt+Ws53bBrVgrqFbfef6kT405U/x
Ep9bBwiA7DlbhXlnJyfCoM09yv/J3QhpnO4cMBvDr6YuKJxhgGV75x7lnzGI8tR4
48CtLuNn22AeR8zawpPZ6/HnDJhSrfeqDMhj9LK6+J7KxlFzPlCBuA4qveWZPf4T
w3ym5vWH/IPG6K70DIWYhF8KgSUdMt3k8ZxgENQaz8nJQbEEFmC8D06tNsmRiBsn
aF8masnwPBIH0AxNR6FcP3WbEghK/NyRGP0fXLPncPQ7y9jkm9hT4nu54sMHljC/
OVkG+KmztJp7klae4YiegG7CWd23WoRI0fAv8+b3Lf++Tw0PbFsAJ9R5o5+nndqv
jRjx2Bi70B8tdW5giidOgWPV+IWgDr4aSqgHbZ/JxqqoBM9mJ/YeB7YR3zrIBN0U
VLjBMcDesVykt1DWnUCSDkxHndbCjYXQZ3xrwfqfQzTAaA60BxZ8WRRIcsi5Q6Ey
gQPofPzDvX4dYJL1T9/dnsvzNXiuagSq/0yaWBbJegF+83sic8e6WnqYeZ2bhhdg
vczjMQmDGcDj62ddhpdVKfQL74t5/YFBwCIKR6gUdemVvG3SrhXVlaaBMqqTwjOv
LNYHpqL9IAAuuLuHvbfZMBKEXMfDAG14IFi1r43ryR5iFZR3wVq2vwMvKE4Q1TIS
LmXra9HX9RecHeOVkLkdgFNya8X0svF96NYJBoV2RobXtba4sxIUr5Wr3n5m94MH
F6cTR05H2d1j9EBTy6bWwuszquoItuD24AGss9o07MAR4zu4H/dpHZVZsiXdud9Y
eFeS+sqeyKQcbosGpTikJsLdqbRn4Xt/04OIgNKs4q6tDeD+W9n7Yk76ROVABWnI
6hh+VytxSiulDnAUTFrNKPsb85YPZa0HuxbLkZsGEMGh2ouxV6NxjoyleGokzK6c
OR6aJ3KyIFXhlhtQLYJeDDKQjt210cgBO6Wyec6Ru/PCD8uzX+TxRA/iEycyuAfN
JaR/lMq1ARm5zVpVMcnLv1cs4irIvwuY/ecvLHsAGoXHHSGmuofqvDjf88WvcNwO
tMRaS81zO7wE9wA/A0DoWBNJqU8MaeusB7q+PEHfrxcZkzsDz+MrVrfR5yEi5N8W
hjdO4Nygv7l1KjaMgP+MXYoveZGkrfAfaAbKYhFi83aiFyrgO6LLzGahRTLWvKfx
aO6hnKkTGFJSeEu4TbhRRKMj4MPoolIKv5hkwUE/FNFsyul3DkXXsZoB3ANxcpqJ
HdciZZON635qQEWN2QEiJq9y1Rt/ALyGWUXq3eoyAWa5fIgHsd+C9h0acKIRTCqP
p9+sl1W/gubGFHlQBYO4rR2gge158+N2p6JqzF02IilC3po6A0RVMMgEBFh5BJRu
7Wr5qqYxWUh4bNvWFaFVf8GFu1Fgj4QTqsXkVPAkqLq2eJVhM4ESA4xm4ajY210M
7qKMjxS19DRX0LJIjXBThBNrPmNriwdKLZZCXXiUp/rgck6+8pcO58VuvxJowJ28
C6KWQKyHb2Gz+IoRCz0jT9SjQRlUar5TmR+nsePwDM1bTk32PSpiDhFcpSq4dJGP
j3SLPD9VDN7BE9EMuwdaHNoufMqHGS25j/4H/j7CuSGwBWC5Nax9l8oHCPPVz5BU
y22nZapUaT5exmIYD8OSl3fiyj5nCPJUX9y9oiOxL3fLJLmPEMzyizEBqGfBcSmu
9vmcIUzL5xEakR6FBTVkPgp4Wx2AUQpmGqBQnNdctzim6FeQztuxMYKxYhSft+gp
lEzXloW1/0JsRRl4c8+XEosvHCBy99A3PzrwI5YV1hbL3tRKBknUfRrBEUy9VkV+
5PUW20AwvUWXyLFCt2ML+19ShdoQR+cw9oEl8Kmt8QCPN3HGYBwnbZUfkRAhlWQQ
t1n0kPDvD2cPFGhOsTbuYkpJNM+ujVLsYaTN2rrE3DM7ShwtMBeNRiEplbIfsnKl
QQhkCJxq7GUy6or3vK87/XArYnSGSdcp5YszjjuxAj4X04+Mvc7nvd6tT4ON1uxp
TfNf/bqQmNzmmVRzjxX2r8JEu7tj8Wcb68n3REXL8P8W1CvrYAW8L/sTJH0czfUo
yeEW8N/n4lzpumIA6a5zN/J0SH1it9hPxYM2XXDHSdA4Y6Ane0XcZPeQZ5Cobx1u
OMM3c7O9b+/4CF+bhcuk2B4ZxBeCmY2Kq5hMs2TRJi4N19Y+JmhUKUefoWtqWpL4
/Gmf+6xSVzclXNFm8yxBohIMfJu7SyiqKXIxkbglPE77egJBvMQfCJQ2BVDxmnyG
47WNo+d0L+c1NqUfCdUgcSVIFAuGH3whMQYHcw6bcg/jvGmX5jZMzA835NNL4qId
2oH1/zpgldqZ777/EJegwwJrcmgKt/hoh08tIAzKjPzytkJaEyxua+X6kJKC27QS
A6oRin1YC9ZJ322eVqgnrGK34b74R5m0X6RJWiaZlxnYgaQ/rSZUGx58rzm7Aw0W
kQZSzn9jmn+aiTxX+dsxyY6hO+i6jDgWORXdfK5EsCnWLRXFVqjsysQB+NKl3q2b
Z9egcyXsYr5A/HnFUCc2UFdrHOPsiNURKd3Ou5ExxAPHHz7GCcf8LIDjQIJz3TqC
lJq0XkuC/3ow/yuTwK2SmfAcGGrj34lOY+EkY1OjXFtTZdrpBE/yWpi637VfUs62
G8kcONPT1OKY4UWvdRIV6FuBHli9oSW6iUSlDMRgYNPSk//fEUeyQq/dN+nuEo0X
EoNioqqfzC2Hg7aq5nnlhtEuOzZJVj5w8pI/nWK2hK+mvDixnWzo3SCtVg/OFG/p
2QlOcG7cXwLaZZYLss7Elw/3tH7IRnVCc7R6rbvYPHBcTj3mK8jkcQ6GKjzxPky7
HlskS0urkJQl6yPiN/NP1CCliTr7jgCiPibRVQ4BJGYBvu6p/NNmcJf4RhySrCmh
zaOqW9UMpr7/fC9+ZgUHoU5dI76DhChH0ME/UivGq1ubPnsk5wWtYeuBrPI8Bo/P
IP8i0blx2REm449XGqj0tSr7QdWZIlT0jR/GEbEqVpX43XNLpoa79M9KmYv5OipQ
8JssCOBDlQL8G1BdX8/UB8Wt5SZ88BVni/FhMmgyi6IvaOslZ623hbNSa3IvMFPk
UDay44zyxZ5TvculVhCsgHcaoHJHHfLTMeg0EiZINP9mjhQYWQzXPuJC3Q9VYJ/o
Nlnj6kKdvVQifwtr57Rh1IQlqPrYKpHpGqjLHOoPArvigQjBZ0ba4+DiKaZv/SYs
g/XYL/cV1+VEdzQgku2GrBBKcOxWGEMFDYireaeB9ldV/BSM/+vwmKdgPqs9f9Mr
evvc31FoQhpoySqpa0mr/Ft/B5ysDGD72aSCxedKxhp3PhdlnVp3mb173cM7BP8P
eENmQ1v02cTIfV+j32vGxJY27hHAc2bbFESrxP1NuJa1RqZrGUQAzgxk6PAHuZOp
woSAvhV9wh4tI/OUWqIh1I35yiHu83q15F2AU76B+xT4PjKnrKhjfUmLBu/UyBMT
a+cq3sVcGmFpcdh0Id7iEslRTx+bbpYFjqQwAokZHjh2mVDEfvE6QCO0bD0VyvAD
iz0E/ke1oQOyISdoMJQcNFS3T2wtukb8AjnJlzx0cBzjHmmb00Kji9iLDt2tIbJD
d1QaOPXxEnKBOzEC9ADz+nzMxnHlslsPh/ZFm+nmIlaUy5t/30BRTzidpqTOqrnu
S/opseMrnp3RJu3QmIvSugAzobCvqiXyl5PgRPlSoyRss1/2uMqMPWvdhzZo2GHI
W5XCOrsZrnu3uZjPUouvOvSFPIrcShOpGuZ12a5cJINRvnxJMrDD//RqU6U5wgu6
083R2Q/ggeUJ30a7zoRz5Xp5JphyYQEQ/9J0F4JJ8k5Gll1YvqH7Snoe6JOeDc49
UezTajKmiiqIERHtQl2fmdwNxh1idBllWoAM6cnG5L4eev4LT7UursIUVi2lFV1G
WPYcofOrbqDOo9L30ndGC8Pl1A5OOtJuTTNHh1nf16w4L280QjtieSI7jHio2GrP
wPjiPJ4l8v5ROuUUzImLUpaEBurTK4GfrdLMz1o1GowVZ6H5YWlMkLfuGcUkNh36
sHOpfOWbRcYz49pLG2ypb7X/wx0WW7B59mrgxvoQ+vTgGmOZ2h3J79n6B7qmVHB4
sfX7FTrFDpjw229peKWw22DqAls6UwOMEHM7HboysGoVu2GfIaHU8y6v768A+yq1
2KNDJcElFLfImUkLDdowx3ofMIP66BTHRDptxIFmTSZXrUY20gqeOTgkzwclvQ0h
pxIVibkV178vk6cXT9uhMB8bhBTwJOiyslZjNtqgKBT+a+iBCsz1IY72aHwLuSHT
jQ/i8UX7QHrSZCEpBmaM6M8FwNy+zZHqMaKEeT9oxFXjc/2BkOrDbi3KJ5FVFzl0
aEHTwwt0Cg8rWGtN28vohdekPg+otnvDxtiGTw4nM/XFadc2OXOcIJ55Gc4SItch
Ku0LHvH04HJHxGgO9atQ6YAFJsWRLDkylhUJ6uWnWH3p/+lAjZPCd+wXE9FMgbIq
EGOzNlUBLsDGlNhAW9VZ3jl1FCDVnHBJAUyqHg+BFeTUki6iBiRkvUbUQO+yltI2
Kd5DNK9xggtisZJBe7XZ6GB1VV4p2Q1tyhGOr3wfLcM9T2OMFiLPmXaKrGHwP74Q
iyYau6LYKOmnDoebddXtSnKpbabPIP0yyU6zYSGA1mCxVlSJm3ftwbWUO2IzzsN9
bQksGhfrALvJ40f9rpPlWDYHxZ+vx8/DWPErseyZ82yXnQraz2RYeVnf6O1FjB/6
5h3lPCyRy0QofAb0uyFkiZygYOZIelKR2J/U+hx3f7t2r2xSD0gy9WXE+5arKsNW
v6DWdIhW2kfiV6VPAeXYS8MCDf344oGiIolSlXdtOVec3YfQpN5br9o56aEGjTIH
I2oR4gtU1rMoukUtsTpgxROtjt4oALpj095VJt3b38wpcgU0IlvO+RQMIuMbtdGV
BeuSF8So6otO3WPGJoPgPKSMVsR2Kyn9O95GEtqPCKp2W6AuSUhXoIwkXXe6bFyi
hKcq74l4f5F2o3A61uOU/AlwWPV7wzkVr+nru7XX/F9PeaLBv35LSy4p70nLTGtk
rHb8rrmPPtXp9t7/olQVdBqplGe2mC7a30xpuxDuaAY1yvK/mxr0SNkAYFvwzvPk
8q2PDcpgZnaRI2MEcOaOHlnZNzy1V6xOG8klXdSiWhhDYQ+F5PyGQTEF0Lw5XlPp
HCOCdJQrFdxhv7Aw/ogwaHUUDXFC67ELjMfELPDZdbm+wyKlQmAILBdcoRJhpemy
9zw7v4ua8xOMAe22dlZWEPtjLwpYTVVeVJcvuz6REXgUybCpnbqOVRG6iizgvC8g
qr8IXUwwY1YM4Is9P+dmcLMy3pA7OKwiXRdJY41jGqGFUAUT3ycMrtlnCw0vTrqL
2Jw+56thVmj3MramxauoKHxXTG/MZLrL5JzwjLfvbSAYf0nztcHm1m+Iz0TeUTyP
lNftnFPArJ8c1AFX1xWx3qSFufJxKnksVoVGfhip9EM1uFYS/PeAIQpdx65ExbuS
oQ9Ie8uvPpuA6qOfiSF3oX+JoA3wzaeiz3VM6dQ6Sc6ZzUzJewvPmWRHK5Z0laYd
xFB8eUfhaEmonQKgvLg3Oj+bmmcjlKbRwIBi2e7HxfGM7qRZI+jV0j/vuO1H2hV4
gw9pRjvn0tvQvUKxj5UqevKjZoCrkiTy02tKyPpNrmSNK3ScgyhShZNp46BlDd61
mTTd20tBOfJpXrdiSakGncYHewynU2OCHqpwPWQXzTVPvd9FuZtpdpvs6WiL//Lf
dT7tTQ8f5xdkiXeRq/rs1pc44DJdm2Vcin4/X4FrVksSPNBAd2GffH7NbXZbYQY4
ZzGiy8VNOz8pTy0siWF2j3QBh79pcrxp9gQExPsQ+Yq0BZlMohc5mV5bsDkoRg02
ghzPqztsALO3tpLZPMEdqk3ug/wFUztAH2dS5JYReFmwN71tEBSshfs6SqAYvP/B
vZJtLl6tqvExGYsQbhiH2krITpuj57U3uzRusKNe9/mzy+uDzDf6B36NgLvFxwR9
5TtqwrJ0KREFAGPuu2ue+Db2gbh6TgQbSb+et8rQpk5nwMdNxXi7RyBL4hMfN9U0
b41uYKNt0oKKRa9+fy1Gu4DZYxHCgXmGTIJOEE0pnWsvOGWu0Jo0h9LXhVQQpXua
4w3VN/SstcWKxOCwpR0APCAWHm9tZ+mF/gcRvQWp3iwOtAiGgzxovE5fC3q/fwTI
nZ2hGmJ5L5GtYbdKCzG0Uxy71PG97vD3K4NFtDKzxYA35rTRtgI4jUT/BCNXOti+
dBG35zOmCVAHgHzIw/b6mFd4ViNdMrTN1tA09qoOnhoPtA4g0RHC+Rpd3Udx9dMX
O+JxLI55lwdJ3X27fMGv9NV60I8hYZH0xJOdzKfgCzUpo2v/tGwS0dJh/BwvlWPv
yJKz4KYPKL/JQzpK9b3O+vvPlgrEreBRUSiObO4hhtq/Cv5mSeBmCliGrTKWy+/T
Xzo/YyLHinTPCN8hIeDYdZfNGAWDGHXynfpgUVJ/hMP8dKBVZ6+sejf6cgDMb1bC
vvk0k5MI+2Exz80xcMyQyxyXaCsqLzaaiwPfxzOAMwlNF0BzauHbuuOFhttl6Vfq
5FbwEhN9anBduhzmb5IaKGr0t4514vgidBn4ixkEKFurk9uvN4KZXIdd5kojZvlQ
WPMU7lfRAZQPNbS0vAFPK/6+qXDM3Su75MP7/AVmm1hfoN7lIvMUbV0BnL19fDUq
kbJuURn5Y6WCiqs0OiNcbLVzWoeZJZxM2eEwZc2dXvHIHkHUyeBdTlfkLZHSX7JK
uosmxsM2RDtAVIIakzFqudEarYu2K7buOnevlWGrTzyO2tV6kUP0bo7gkEPt6lz4
hY2Q85VoJu3k6QCbzkqZwAMQZlNM0xFxOgGD9bxQ6ApN5iqsMT6YI0qeDSMnjdLS
FMC1mLBKgAAmtMQPUpzwuDWHOWJN9E7pI6aQR87bzU6AgFFCvH7C4VGgZ6iuUZDy
Gh5PxT4uX5DzbRDZEXsr2nQPV/Q2O1aMUBKlOXHRSESqZY3OnU8N8VDD7s9TlOFc
VJdyJ2gv0Xmx0hJVHverKgIj7P2NauBKCQOc49WCTYhEJ3wVWQJWA2GJRXO/058t
CM4JK/SL1/45HzKbqZimL/Q3ttkEjfhKdG5HxpsZWbeqsRH0atDGOwvHFof2g6tH
sFsdDB1oHDF+bFiCcxq5a50REAe5oR2v2uVjVFMjgmeapWw0+KpxTkktcZJiFi/N
5MVPjSZZ3WPjNKIVj9cg0ItnfkYx9o0///xeuW/Mrfl+5FDje7gdaordj2X6BAzN
FDkMf65IUJ3GsllmVhXF2TpMgCCpvu5hu6ktjsWzO4+lNQabbqkQmCodLAHz+DSy
aYjWq+H3/1ozGhYB8f6T10b7ihwGXbkF4/hTNVAHWnlWaUIurlZcf7b0AL9zjf4P
KRJ+TRt/8JEJR/YKyEq7FVPxWjr5DilGya5B1Fnfv5vPJYJDaGXezc1hpxmivXTm
bRxM/VhnhQzVmB8qvY09mYgxDAKWVDOicqRLfB3S3B9LlB4/aXNwIwVLnKFnp3fn
bLV4zQ0F+VJjzmnvQ73+4U0gsAWjQ1z7p7wdcyVQJP8F8V3RC309LOYs9twMqxk2
WnTj6qzqdz8/1i+KQBJ/YVMse7RKg0sdUy+Q/y4X1nMt4FzbJ6P+I+/Nc2R069E0
UoxFkcKdY4Il+EgEJ7FnLASGcD4COKLmASm9KKftUdUQfow0j+oMPX4MwKXkeg4S
7At/e2G9EKB8EYhrh0tRKq0njj4n3ADwkdgjdDEp3ZYpKHBqTesl1jnhfMbJyQcw
V8oBBjre+EjT0lvKeWSNPZMFuTe4QCO6o1Z5gjTUavvCO6RVxvJuL0Kf2wgzv23t
nUh8eYRXp5oE6IeG/O9+kxlQ2IQsyULfo0g5H3vJ8SWYnOXc/j3nr1HsWruq1gwm
D7IhUvO58VM3ghNLyfiZTK0PlUjkiTnHpb0LaWyI2/9WQT/xSP17NU6IAbzhsb1y
GZO1REmpSguBOFgbQ55sGA0OMix4ixNcB5ix4G/eRV4/RYF4o5LnzMud9G5/IOC1
M+rLBfvLfgVGcXWxOdE4xEoWXbSli7mflxC7Ys3JSL9thHZe09BbAr4gZ+wxZsFS
pI65q6eP7e7CxO/fmYD3hokVKxw4n5n8V13cYzWlLgVh2LQ3e6Elis5jjRxj4c/f
oq/zUc4MXq/O8y7ZSL8IzZtXdN7UwmQfLQWKS6G/WLohHMCzLCK26h+HME9EX8Ej
yDXqlJ5hle+D9Lvj6osaZQrR5ZWG37mrQ0us+rptq8Pa9cAP7DItvqqNvgWLYT+r
+UCiyX5jMMx1+Tp6573IMpoLuea/4LbyAIv2cviPVYr51/H6LsgNJS/A856Ji1NN
HOhLBd2M8j9l2HIoQu/35yFbH0Z4SDNznX8RQpw4h175Q69xab7OffbLveICKAnw
1U1QekoLeoMDmB27vgLrfv+pqo2ihD4T9XpYsWfYAfbo3jchKBe3rpik1VNkvbYR
09ySas4dzlpV+dA93VM3NuIYcm+4SKB9gJxZAVfaDEz0AYhxre4iLCKUhut/m6Hh
csMoJpKIT1SZnYGOW8FqUza5vNOsc3zcIN/fu7iFP/T82U3zL6TR/zdOSUX1mtWE
GjtoUjV3quBHz49iyy0O368q+KXAotp/C6r/wvStkg348jmVDTmqEKq8+zrIahhA
V8Ur9ojn6QtS+rkLcaAKL0/VZqs7eCYq1U8hV5h1YaFJ5vVK1SulgRQpdk9F9hfT
PK0Xy2RqDM+FtjuWP66oDDohCDmKJMsJe5jUT31cVTTYID7UaSzGB3PXzrFHsNaw
Pw3f8AhwT7xNgXhUeHW+l7iLSTvvaj8QnyOnUF2dD573d402TJafwmQkfwb6p/ZC
TBXJuNJy1Zqikw8wMq6n5B4azs7ILmTUsuokMc3whIwdDOMC7gA5M66gcUbwBtMy
p+k2JpsviVRRsW7kHYkCmbTj6f2x67ojQ7SAZeTGA23g8RWKN93HzdlLni4GNq2M
FID+KBKkUlCP7N+gqZvow5wDq+CH/7Jb3SGLKvpah5rJbO0PgbSrOsarH5MfJq4z
jFjni0SEUmpR0SQhw5wCsWoZYv1d9ReoW0o2f8GQ3YxND9adKIKwIhHToNd4mgzj
Ct8z/7+8SW/JqRRDwOzsBo2xSWVfy+xYxgyvq/pF/ob76jYQeCCdZ+A5stdhW/dJ
jPJXxf1xmwUwQFj+nCcj8JCsujzy8Wvryh6cnf6bTp2d80Y8mHCI1kwW6bRkUq+f
th/Fd5d4fsenpiBe1qyHKx+Duq4d/3VomUh8Yn6tnGN//aA62GvLK1DOzcAJDo0M
2GidZ+Gf2cvTzauqzecnJVsPxExXsabjNx/LSfkqPlP05cDznnzid9IzEEkY6h/K
ZgfwT3upAkY6IEDWjhgxwSmVhAzJeiBr+5wNah+aVsyNfxlSCQZj3N/5Z22x4eqm
cwqyh5Tw5mhCG78SsQplHEq7Q7aeNY1DPvoLfesjF6LcE+23hnZdsBSJuxRUXTbI
B4lO8oyAznyiOvJToskmO4+NA6txQEPR1ABtRs17n/v9KmAQg+LgBUtLAbwc7+yC
V7rj7cAWiPvZcofvTLYx1Ww9gPAXg8Vhkylw+98A+e8mhFe2/wCwIxnN4OWS1hX8
Jr6uCDf7GomogGVkpaZq46an257R6auOUDfsiFf4g9hs/ehfe5YsV73qndqXM+r1
JOiWBHccXPwaMIlvkDZV3hxccw+nNuwZ5XOqsDSnfrZ1nYSx8gHHSphlW+eFhkmI
+FX2VQCuJGqk/6YsAdLr3+NntUrZQ4XCLcZMURRglVc71aQqXGUKR5oqYYDwkTG3
bDGVkt+nTVK6hTBdZ475zB3Ou8g9fRPE/eDyOorlX6mBpsCICH7chnwk/UADBr6O
NecBWDTY0ZfxxpfiB/sxVgAVo979qvZM+eWwqX8W0PtO8YoxIujwBtnznGlLSbJ/
p4fZlKADvz/BytcjTTOa1ughcaQlKu3jM34uPwEy88H2SLt1hTTrrhf7+ehFT6iO
mW/bjoo8ieRe03/Z9SEEHEkLjiOxjEvy3sH31aywjzMfikDhGo8FHHIj7uvMestz
a93FY9NMtjG7l59EL2+RzDk5gaJPl3ioSQHtMlWBMHP3nhwKXi5Vir7ux1m1IJSE
JLcbxnDVMDbTWgLdpNgSLNi0FHNyHO/21A4luiESK8WHXrp3KxQMn2sF4JVw43uj
5lecnqrgKxCwXfxeMayCJNKBrF9rd4TWDS7GCfpMEXDpg4myZrDPxO4pi8PkH1g2
uXyBr8RZf4uBzZFr+FbLmUQQpM0FAK6odceWkBUVBm3Mm4AyioHsv4WDImHnDrKI
GE836aHerKjPz181N28IhLXpZ1R6lrEauVECphUc20iA8sn/9ixNS+GGSF56pAK9
hxndTB04ewHVGRNt913zrfZm1iZfAEv1BnVE3sNKNOcXPZJLdhXDBrAZe7b2PT1W
aspIo4D5f7XO8XQwIW/BPa5X7tkLS7azl5KhSmJVG7CUckpHhuB/ZlXnz4Xy2/mv
p4Kv8CakPNHW3o5Bx4Wsq8UI5z3yZFOqgYqEJo1X/fXdPKEVSFEXOaDdJYG29SIv
UcfXroD8uzKzJNcHZ6vVNxTBgXOxhINHQ15U2u+gvs3ATq+WjqaRtvLAErg2Zdc7
AbfYFMiudQ97nW+3n/STsZjhOti+h9iiLvfqWAIrspxX9O96sodaKpmSG+4KE1OY
3JdfuNYENyejn12/XfhZqCGYmH1ctbdYDAZOZ1kgMliIHZA6j49GHxzKI9IfVOF5
qLVpC+O3SgfPTjCIO7qdSmm/nVG/JLNB75XA2CDAGwvcAEXbiAEIwTqGE+XALxAk
//kWiKWsLBe488sApWDd7L6fPFGWN+PjNClcrhu1YNZ6vCPD7TFGMjI0HRFCTJN7
+z2hFQp4onnz8/5Ou3ZHYB7tCLHlUzUf7AAL+/tixgQuMvgA8CmK14uU2Ypcylsv
An+ur/A/bjM3pY8Wn+FL+HR149yPihwxJvPH1OWsfoEJKjerAwWcmzXAFchr/ya6
R2/YQ0ISIuc24SgBa1YvxotbzNsNgKu0ZaasoC45EHJzxdkKrqM/FQK01aDF6lXS
mS7bHoUzheg9+/vFx6z7ja2uJ+YnXz1Q0hXh0HmqM9iVxYutDPG9x0FuAckqq7Cr
5fEY8bP/IBfSA1/uZnozittXYt/tt6UqSYlA2hZW3EmtZMkc1footXlTmv7obzvt
IrpvoE/wMr7fl7kWq3wEj5sUGaaDRvN8sCGLauEd0ND0PbJmk8ygkkEJha75E9+J
OAYNN02GHPGzclG50OzE6GUOk1R6kdJEMx6q1VJZup3u+kdpAnxCW/mTUJmjLzqO
lZRlHYQ5aMWkYJVriU4NTHN1qhE456Cbf4zmzWUUa6R3Ae/kdxxMAL/3f6UOiLDd
7XkVXar01nuFQu0KYPq/kvM5vIRIhmNh93PL8QSpmvq4oy8cvLQwyCMJe2f1WjY6
xUeKTuwveLpcJF39T9+y/PoX8BEv3PEI56p5m5ctn0BrIi59Yy5LDTpGM+JfC0O8
+5NFKQ0+QmaVMayr1HI/iYLCd9wAFt4JSkTTAa6biLE6AkvqH/pV8NwSsZ/uSIUH
ELdY5AwGyTwDDN4nG3cUS0MRQcSoiLnYjh5tzbQpfiKFcH8L8VmsNNVuuFoRyVXh
gE/u587H7zi0UEVG4TSR3+3JW7BDd7vw0jglW0ScPck5SgL+akzrqlgqC30A6mmO
Gwc4lT72/wbFN7HWr4snGL8XZhwSCJEER8mz/omKhl27vXX6mOJ+CL9hhXjtEKvW
ZgqVJdUUAJ2QA7kLLjhwYR6LXj9kB17z5zZefd7Nx9lr/o06eYxZkdpc+9DpdE12
66/13RCsq2zl67pEZ2W3Vr//vnlLg3SM8FbeUQrlfPInHeweuJRvzNZGmxpBZN2Y
ZfdwjmkfhAudetjjji+Wi9ioQl0A6YO37mYzmNkhqXfgtxN5qQ0jHtrDz+34FK4u
HNVJN24au6N1orVObbVt1fnogP0PEAsIjT2NwcMYWECJMyVzDvoLFESjYl1pLvcX
hvMuC0YZphODj+zjzLbZoogJQATXbsXoR6LdnHqQGLvvdvtfT/C08uT7cDl1BO+l
jQXsL7MfyLcvcHpSjINUHUaVOyvuOfrx9vDtkjxacFmWuonOx/HYVhSL7NonGKKs
thYR3lRGoYvcVBdmxniY093d6EFM6QTM9LK0oaQjSQEcG5saCB117uIxsqCTkchA
OyrQSgafGMOAyyo98oiHtebOmrFaMJ9ZAV//3rprE0c95wjqKmyqyyGrm0tyQ8x8
DAFhmUE53BGcB83wsXJC2nW+ojy6/z+LSxOLokxFw6uLXKgIDNN440Ocx152HUUX
L4guhFjpieeMncvzACeu+8tg+c1pgmPhefkehfphAuWKHM0uA25M7G/SpAvBQxa/
IIf42p5eRZsv2T15pG4QBr78Zx111a90XNfF5SVnqZVAp+cdSNIsQ6Bl84wJoFf5
1wD5AJ/GHF17ktpAWlim0XivpwzMirhiLeOg5KkxpmzbSq77QmUYbAsyHy+M0G3/
SXf+Cn2e/PXpZfhDRbyyc/FIj3RmQqwJnioVeml+whBCunNyS2h8ZyrzGhXLy49h
2hr8lLwXokBLeJHfOVTakKEzTYt0aYckL0gw7t3gMECqDx4uvdNE+tr825BkXPdY
dUYOwmFLM3nUf6sIVlAavguYlW6K0+E9n/ze0FyD/SkOKpLXe0kFxR1aZtxV36oh
yuu5csfNLqxW46Z3C8QwRQOxNqM5BWa0aHznEH26aLmOkAtocxIfJrxuvcqa5trs
BSH392fvYuwngBZVLc8AeIc8yTOaGQagQI4xEDhnPQzKmOVnMlQV0cIZoco/R/3r
QOnz182c0HLSX9aCPkE/DWCSyg5GcSCY8uf06HU8ymQC2Y2LB6tRgvmATCkUXMHF
bCMsykKAcPFRS0DMFQ6u9B4yHmA/PnqtUb5PQP1Hndkt7+gp2TwKjXmBcJ0SsN6i
xIr4TmlmiYa2ZjAv3cdMeupmnccK4GxWvlvqk+H60OwIj8WljAeL3VfaCQ1VL0N4
4mDRZpekkJy2rYodcVzvCJs/izIQvE76Lb6Wx4MtcVdmx+iN7PLgpo1jmCJ+cWML
7E5kVyxP0tCQZy/iVnKa3WnRGbbh7rzJXuM+IgZ2PHZIt2IkvIM8310LoBQ8Zrs8
Erxu3nIHkco+PJEBnS6C4wklgx5Zasrh6o532WWtdKv1T2HwFWeBcgUNhg6lLiS0
XqnTCCQMXotWjodRoQV+c2F23D1uEjjOfxKNXThJVTm44C6EISwOFS2Tctl9jMwn
P8RAPCVJYT0J4F1t02Lys6wxeb877+ekfeYRqF861GcqBihmgWgFgmByc71mJhBS
qqmjwcmF8l0cbaXJhvFG2Mv16RVAJzTTzdQGn47vuQEWuckOBwGxvadtRyGDfn1W
B3LglyEI95IftvguIJ83Q9kJ3DZ/xRF9ZYNgnHNOSUXOxBS7KkQE07YTBIaRg4xK
hGOKRGChk9p17Vuqf26TcELrAZIx2Qv8fXpi/UFo8Lg7+M5HkFwKDMwBlJ1CFsNu
OBdhwqnmygVnCtY6XZrl/OudfOcwY/Vo2aaiFaj3AX4zw048qB/GmvixKpe9nirI
bkM+r33VlFXVfd0co/G6a5H1Cfq3ivp4GfRPtkIFELppwZRewxKeguNkQaoxS1l0
3rppA5grBsKAfjpld8z6vrToK1If/N1xrWiLVqNhqa1dnN1/PayMeYXh8yC4Iu88
Lu1hNHoCxPCf+jpWe7GtCvd01d5XIiH4jSX8GbpNkZzdX3dFxIjVzJ0Q/fjFDhl1
8KKc630gd4FJogdFk717/zL7Rf5+ZI97YLRwyMTaTMN+a5Uty3/H64SJtDxOZE2V
6YIS9z2NSkFDD/wkeNjQ/RnpAuUkswlSGTJUehUUzV2At33ow1N9tkC3xJc49ik7
M5ywSKTuDpWQeUVtrwLc6sSDoYR7S+MXd0PqRHdPglUWO0eeyH5N6YBzhHSjJBW7
ro8VmD89j0GBGuxO5qWdSRHQQEIxEOGbbNzx29z/e8F07z6UiH567kq4TBwMbAIN
pLCTJL0zXTbn9FSTq0Y79N4APti+u/OzYla0auzqDHvFFVLBIH3I76MT/PLLhmoO
Dma1H2fM6dQaGn3+Pnpa8UZEMWk+xGR687cuHcxZOMpkwBghUvcUaB99wesikxzY
qdfi3425qS0BvyQS2laGvalyqri3Yntqv7UrpZLcyy3xbFGkgSjZTgls9mVRZq26
IVyljZy2OqbMbuoa6eY4GtzEqOp/cthrQDRH3/Tfk43RQxlaLNyfH0JZG/DTwdCp
PBh/oFmXrFOz8Yuaj1RxaIpjKrUS948qvAHNzDezgS7RHYKIN0psMiOuEmDnBbZd
MI1iRd3b6Q2+vbyOT78NhjUwsAWeGEigLQ6ZNLv1rhkT74aEUhpsHrzzRh1imBrP
7RVYMn36xMQxM8lBPTGOZ63mDieXbRK+YhEAKlWgGhLIQdKhbliyYMIq5XsQYtRj
KIor/uPg7OiLHVqLooIMrevFreQ7Gi9LeYQGiWbDcs+eASZoPasyU+3suFfgOsY5
Huw+L8GXi52uu9Fg8WHGC65GGDey+fJ6P94KlEjfe+tK/rRgfA+Ot2dFUkld3kwY
66NqPnApheey580Qmf8DBCbayLAPaW2lfegL0qTPmLEZpRGC/60mrg7BMdPEuviA
ecYUCiSn++/C12txEDqMlgELWdRepIVfSwjwdz0UK4soljoKfjgvzYwnaKkw20AM
YXUmrpPmz3o20FsAIG8sMoQhhAYr4n0Qrh/1faOz0KylqHCEFcTL7yw1LgZdjBd+
3db4+R1uqlkPTX31NL199bTivRIXa48QbwZ0qufqmorZExKfWLAhE7y+8cORP78U
0PAQ7jrT6ItNN6DUZShMMCToNWKDXUWiaAhasQb4K6qtIJi8r2BY3Ns9/KPVEj6g
TwBj9mZYGJJVrmvhgzvMsbZG+qyLtzzizGTx+TeTaYP2bfE29OvwNy10A5uC/z0t
BQekOQTL5OmWOimA9xjIUaaVaB/GW7X1a7D1xtl3Zfve1aoQqg3EIFn/nl3lo863
yDmEq1EVFeGPmkV9aX23lvckiEa7fR7c6ocfYwo3NSZ7IC1+0WUrdMOpIQPX+0yT
ZxGlX5Q/Vo+wpLNQ6fuMdw2412E2TNb0WmUNcvXLrbGF+9evLgYS/g0bEpdNvBwy
uPpsdKOyDCjhKOr9/1yIzbJe7jIpBi7HlzabXLB6BmnzsCMgxFBT8xMdgmJWfxry
tz6Kc3JRz6/unVWR7KNclIsGJIyZnUSPX5ZvqlOAZ7oV8+fGvrFlTVe3Du8dgGAN
drfhttk623gGhEfSnWZvjwVyzyDMIOl0sy8TfG9PCY090A2TtQ9QctwVtK27TGQJ
Gto3zXz6Duqe/3ptonPhMxPUXs6K4LS3+PB4kMYpqLvqjv/1+OvMVPz0jexOiWTe
mK/kU2WC67MEUfZ9w6gl1sWcF0P/gRtvfvK0Ses7B629N0fS4JQQ/dMzoE46XzHv
XgBWlumFJtLP20Aoc4UNmSsxr54HbUZd4xFo12sU4CYwtu/iLUZ6/XJSS6ck+BNs
2rmc96SLbzHNRHQJkWDbgvjlyCeqs+ti5ePfb9OKoQ4tzYoyeVLr7w3w/3qezOk4
9F1qgI51LIiBcyE/Dv01kNmP/nDVR07XCUAq+8hoFgRPEZwEW7DCblK+b4IGRO6d
nhPIW8qE8YiHH4iPQemidgHOZ/KA0fvSllxbQX4xdFP2REDamZvwTb+BK7zquGB5
nXC+EIMv8qZ9i7GLLUtTgyyQsQgTmXby4WYy4vZ+jr1YVmu9SutnN9MteiGfMROe
PkkwsDeFv/DnylhDGK5JHV2YrGryCMg4CYNIvasBGBPvHJaXS7SBRNJsKyT+dDPi
RPPaSdLH3BgPf29mDOJvYgVKYnZNqv1TLNffnHtLG4fD+/VjdDtjz/J8B7YK658U
VA4IgL/0+H/69Gf4RAcwH83n2suvWvRtm4VLJFPjndLXqisgaSmX9rnY9EqFvDnT
hiMK4RgbrLSzB8xP+enLLgWlCDA5XJ83NRFAsu1/opQWtdBoFlL41klTwxr7LBoj
7bozD/7vXNwUF5xz1//77IH6TzsYpAD6q+ZZ9bYKBWpiSIDsNI/5548KeFyV2Ru2
0bZOeOoQBw4RIFvSafLufu70pzmRa2U+SelLmNj6ETmT8ppIeVtCXWpFw7ZDHvQG
VkJgdMeTFsvf/ac1yLHiS42XtpzHTW5cPKnUX4dUIbAUYWvFujI0svFZdSbHVN/W
iCvK3PT7wzJUrKbWPGZCOAsnOAyvpNh8RVDuhBUioRWbKWduP8HO6ab1l9JsNBYk
qz7y7z1TXiuNNU9Xc1ldg+p2+Gcs3U62wA44lNEb871b5ZK3VecN7JvjrfclJem3
666UfXzkvzDtX77iJOOVDyUSfgiM/1uO474PayYuYIGFLwKXz6DrMzGi7hzSGe62
uYOHygNqRBSRhQekgtaBYE5sbLNriRwGz7JD8Px8SSddTgQSxFGelODSpflZEnK5
mmmWizWIUSxInA7kPt2L0AheOt4Qpoi7VLcahBizSpJGk1el5HACxFNNF0ZpaY4F
ac41PUBkX49J6RQRAqNfqB1dVtDKA4S5cBnk3/vng+xqL2pCLVXJF/DTuqWKIib+
UkZKdkARj0sdUGCaQ/gqOV9B7XxsCYgiopJnXBRXfwFscdgxCr/h0XJ5pWz+NczV
KIWFVVgl68EMWHg+MPuI3jiB21ng4B0YukSF6y6/WC+CDc+GesVkfxIJWFoAADao
s6On3VGSfj6lNTv+Rj1PcizO8Jiyg0dDKeenGd39CgILYCz3SZe0M/fPov7gLLCE
1FIPBp9JZSfPE4fJ4UYg6SZS8kqRWTkUzYqJM71ubmSI+tuQ8Ax0+iyRBS0GqY2w
R+1CVyZL7WTguHApEQ4QKop9mfz6QUhrXx9sdiMHx5erKRovuIqX7ZTEq3D95NvN
PeaF00Pm2bvFVQcUo+yk1g6RWfw2Q/zC6UUnze2Qq3TGeqAJMI1DDH9Y3hvhpqHS
G7LmoPKWizkNettyVMo+0/x4+9VnsKFbvkE8M6cTmunsHuNMBrUVy2yiyrl1oVvf
Y7quHJ63n4qYmJ22i5Ly51wSMvehjLcMKp9pKUmZmxQdpcqJoTmJih+RmGG1SLaX
/K27L2PV1aJ7hfM9P2y3c9tX1uIVNDpEn4du0a/QiEPYsNHw8sqTYC7Axp3xc+mg
Dsjvr02M4Q7jPk6DYi3Kws/WPY15KKj3MRgBU2gU+dCqsyvOWiD+INkRQPrJhKOu
dS/Sdc+zZ0HEgnTQVcTxPFTRk2wyT0kZLjUQtdzCYVlnrQLHaOEhUKARcGkrRdFv
6qcA4Pu+ZxXzGOWBrJxH668ocEDdcNlnla/dy0fFBdM/BXf0tYhcn1ccE/fCtiJd
NeLMDzFo1J1Uj1ERplSWK5eK/xgzzV3/FTEJehWD6hsCNB/4qLiUcgg5dMY7Yq71
1YoJj1DpF4cTAHVbiICl63hvJwHdQetVFGQ7vNkZe0nmiwST7rdwUVyGb9P5uTHT
x+VHqky0c0SwGZoj5wEsFkbfQqLSPr4ru5EAqcgttvUfPitoUTSZivDFd4jhSivc
IKvXxHqpNrx3nLfnzwUwgdwDNLRZDMxIFL2R8Knbeior/4POzeySAmRVgQSg4KGp
YLZmwOOcqRhb44L/IrFT1cD3DNMN1mP8iiBMAa09u8GzaOAmKCk2rH06dCovkLdc
JWJUxLOjZ1/kohv05YN2BvrACovlrpi8jJGwh/GhqneusGXAnfV4ylo213U7P8J4
NPHFCdTpagddS4tlZh2v8Z2bHK+Wt2FTw5qwg8qaRrtAQduhNwBe2IU5UJr4UeVs
vgO0jwleR0auWtspCQro31l5KzJYdYNI1i1ifhrI2PDFZP7yx15teaG07ulng9QH
K4SVwW+eG69hGhyqStuynkMERM/LHZQWmVUU09mv5vQCttTs1BgCRZBXdycALqcF
pkgpO9aNjLATT1G4qvQnlxX3leuLjyDoM6UzPpjD7ZpmwHS3QUGZNAN8B4Rz/6A7
fvyB64N2c5PMb3em3sLhTYP8x2WSbbnTryRev8IiaP8frRUS/bO9MYkpXwzky0tP
5/XsJrpM7KGPahCK9O5WfDPFRhc6bg6gHzWieHHIVf9jMxydUZQHqdfF3IF8QNpu
p6vgx+XZUiP4nPJddunF4pT7HSO1/zLmXHGsJbaU9gYtOPHOkeL9eBNinPmCNurT
p2IF0mhrYxq53DJGn9my+tIujIRgfKvp7g89ewqDl/KpPWebpP28zf0wz6eBggcs
GpSz0Dc5dLHImDfKKdmvyaX7jgQcd3W2N3IG7cO17IcT7YQ223UwaMA7Cn5HNYG9
V69kvT99rsWeDsWby+rxA4Z+N1JBTY59oJbYikJgdWRb0+lU+lEzibrjvzTX7bPa
dhXpK327WQVLd6SsvPPJlCYfpSTXCscyfAjGuv4efZXstY2unzBcT4MwLIiTihbg
fjpxmTcf+nrJ09i9YbfO70ihMjXsf0Sfikq7FFs70j+OKFUoMsD8YOA/0OeoC3vn
GpVb4FylCTmh7OhiSZfAV7pRWePVJ1scV13dIi8QBvZOos5KWpX0qhdp8CLj0g8i
qDhU87geaGK4GArgwEaGYeoTvwSD84fUEJL0uxOMYjw4NrgoUo8PW75UbNBHP+S5
TQogUa8ufJCykyTHnfjWqyIvQOgh5nvcLTeDhCqFxOZ9dRFZAU5Up5N/O/qM2fGH
2F5R9axpF7UKrw/FNNbCFJfyh+r3tqILWeYpEpCJJpxwz5o5+9JFnOE9/O6Dcysb
xv5HVe6i3tlSouXGpKN6ENWqnFWdbJfhtprNL/cGZBEh4MedazWm0s7gGjZ4s1tF
OVJSt/cHkYfr8zM9NElgSGMjQp80dykL+umGN2WAuqJV/RaZZpQnn1w0kP+EGJNC
zPs7BZ/E9ElgjDR+dTsPpjBOaamQQp3Jq7c/48OdBj2EDjL+urpcTrVUfGloJMHq
HpAIaW5WAT5JYT1+NKasIom7XfqveUexAYmX1sZL40WoxsTi9iqmQfiPovKKnD03
jtH//IJkeNO+Zv6im7X8ogXynlx5mTF66H70WW6FAGj+BfyvpLB4xu86T3Ch85IY
Mt3ApPyHOPBFqhHmO7Wf1mLbjIaTXil4pMoPM/hTV6UFEyK5ssyF+JnftkE1ctqk
oIPqB83gOiIyAj6GyF2ABhWafNeJswuukrxBZSatv85MgDUfbyos4zcTqFnVWi22
DCTQGFOq23e7TrUMQc/2OillcvU98oClePpnXCWWwGlMK4/yX0YEZMVZlyEk+wSo
FhlhOG78xKtvm10/0PMnd4zL/Vt5wRJrlaEPhZPOQ/6J14+StF7SZQrZRq6PSi1A
XmtBr43qgovxMCjKCw37b8AiNc0Dbah1fh1oFR7tDGfKYRzt61jDuvTDfVz33w3a
pMdDFEw6CwkqsJtVqDZ5nYNGdv7y0AbJ9pCLotSF8cJOgh70hnCJ8ufV3ntvWeJv
lnbv6gE+7ppN1QTrbViRchwDc576VcgKnygvBfGMQFVeJaU/pjry8YjhCKovpsqW
SGgYXasfOl48RnuiBCjRvdGoKOuxH1kaL7LC8IV1VCi01QUog7/9S+axsN8/Jte3
L7PUC21QtV+m8Fkgetap27WA904HdjrECOkCGf0TaLAbrHjNVoqcvWAe7DKvIRto
58+9f+cnqYYKm8LVUtLysR/KPhK5qcShyNPof9rQCqL6adArjCfdNPYfWdWei++J
t5vDoPPPxaXAJZPHeCGb+nWWx9BWnjlQhY91UPTv3haEQb3PGExciX4lFNtmwhBn
Y9R5nthCPuCQzkBIn3gFynZxxGxROPNQAbSxzqikyUQanGqKyo1W8GAC2XqFfiv5
WwYLoBsOBAeZIZAnv3RiEY1edUZ4cpsOQny60uQbLpGDgc2RMRHnJF7w5TXBgw23
Xf3f6v/iimekeaQ94vkByndSwLo7cjuCSeH4jP2+cvc/JwZhZ3VklfE/g6m7Zski
rxD7k6jcVeMexY7PjYkr68t1MR+vzRceQ6lrTMXkrIYo8A1iinmrrF/s9GjQZVSE
Jiry0oQ2EazEiIwrXmqMQpfF8TRol1Ac+d4JHusuvBMWH4ZpAE3fJ00CHzdvAgBS
o1K/aqJKW7i3DJWVyezKSqUD+XYDtaB/1qlIf2eKxYRJZyBGB5JRttm8Ayd6UDnT
eoDb5BUhry8HxMbP4jwy3p+V3nhvvgm7uVDgtiSLY4Db+YOJfEgTE3cPdT3AWEL9
rvdbI9Nk6QvVJbd7WBhGoTLfC6CZHy+iICWsqm3RzdM9UvXk9XhYq/xZPLsjzEWv
8Twz8DnBHWRweGzfKtyZXx3+H1wvgyk55vxfYpio7m1Rn32WToO0vJZMboYVa0C8
nVJvIp0SYiD6gDAeY85RkcEW742BN2yvkZZqUnzSGKQRv8gDD8nGmEUJyyuB7/S8
2qyt6sJoMuB7hNaH5NbB2QhbhdKzqkmZxPbZNopLvtfWSmWMwArXz/WDbtm0KJhx
/7ZJ3URGrp4U/cpy7NgjCwBx2+ZhVW3+Y3IJVG1/6c54MqogcvCW/YHkViBnG3Xp
ZYxlZDBjmyLjcwZA6CcFgxprrz35UGS4C3+DUKyDdKOsXgNwfXlhPHqLJjCTFkWk
wXspUcKmhBcZY3r6U7QEJ3iguPQ2GwfhySF43tP7QLS8iWXLcDIVE9fLhLyaGW6g
32XV4z99/Kiv2QFD6a/kRrjNV7yaT1tQerrH+WyqxK4c1JxdaHWVXbaHcle7xQ8O
Ni684a0a4HHNR74DOXIILV/UJSqPeS6EfTBPg2vVfSOy2TAMqxrv92jblibWXqyq
KdMDAtTQJLyrT34S9qK4qQvo8SZBIie/0GUSs/0HEThNwtUSn3kb34HgdrL8I7nP
ILNTIamg99iQKtHFZ6AlHANgz0SkERhM/8SSP5JbId8UlKEINsYB2yIB0J+molao
Zl8fw0GLnGNAVZKr8SFcPXemk4j/UwjLrK+qPDxHDQL9jqpFbflGQMnyraKQbWGp
nXpP/1FqISG3u39xLxWA2ue/lVZ3iaKMebqJq8YYk4owOzgpHZn/C4ZPsQII5eG4
YFAW/uUR5+ynjxTrzAVu4G6oJhxxImyJEWZ7T/gwMDdJ24mdPzzprHfh/1P2HB65
+sNR27nnZGVOlAPNGJyxnCj77XVy+4i+hVv9VxHaTpIeeHA+4BV55pabU8lcBL8x
knLW/GnvxAVP6X6VwGdJixcIGh0fQl/zRs7tRTAoTQzc4YmkWQl3wnCqoUbgX4TJ
7/eH1G1U0EPUGMiEthuUtMJKH2Wd2NIWeVO8/WSu+H4sIQJkq++9ZIiCvGywlGDr
iP2uOZFpXVkmJ/ANYCdMdgN1eergsTK0gAC3ptMNFQ1PXrW1TrkssEYINKjKDgnO
InkJd+KJCG3IaNdU9h1i5+m+gXcSNoH1Qiwz8hjwt7h9aIjueeJXBFA5sK8mvCTJ
3vQgBhyp6n0k+bADvpmnqeG2nPiwn6tNVcopaj8XLb3neuA6MuGs06S1fdmIn5dU
bJ80OolShLOQJk/kijdgO4iB8e3llHFcc2vOKV6c9PPalKBG+U2xuHNw9zw4EY+q
7CgQL5VSGHJBJY31rl7JFVDTHjAfoOzC3lVwPNuLebamG0/Hx2ow3VN6GWZLeN7i
oiaNsQ9ivATp7qPdsTwpgyAGlrVaAvjal3I8sxcCBmeEY7bTu8uoIe7M7a+6PQAD
OFKjriMlwWD8B/bFTArCY9MEAeyNCauhIvoEvcFwTHdngW55PS2ML0Sf91AaFTLK
Q9dxZZu61M2zJMUIcdUcQf7+NPRbRKJA0v2ziWGyN5h+48lSd3NhjTjTSXeenYtI
hk5endLF1Acd8BG02aZFFG4bJS57MlNKR73s8aXMiD74+n0y94k7KqYy4Bis89oR
jX+1iug6rzDt/v0BBhQ9G48Rm36eK7McEepIjtSNw/ahk23arfyMDYUNejC0OHBm
cTbgtcWQMpN0Ps9FKAPU5MGtA3+zWhdcFvfwM9/frkXlpWf2u30GXxiR4KCnu9jT
1fLt76RIlUgOo+JcHO/AuSIT14U9xN+hFC8zH8ZxUCn8z2E9c/ZMky1gey7/aw1m
XOaPJYc2gY839PMm0umoF2zWQ3/cr63JhzDrzapt0up48Kw0q08MJbnpL7gDcIjv
YIi1z1zJRSoDi6Gy4cgNImxcC8Q1Via0yJAYJoa3l1ZVKIhmBmwRFKhHe/zRfe4j
OuphsRSQkTavyrxLaKEvMOD6jqFzeG4HuG2CYdyRI9P7N+FGXJ+BcIPScIQkTcmA
MAWR5Lmax0vOOyGICpuzWk7qUWOo4UurqB/Rar/YWzStkRVEr2iu/uuXtntnCOJ+
jnT+3XyceU1Lp1UXhCk+DmhgCfv6zJNM539y46bMvtqili8hTLqlbx1w9C7HeLOX
9M8IVlsHdr67sgR/juhIvq5uPjCytWAsb5qzNYG6FPKhOqJ4nErTIK/seAlL3mRs
4zJhfo+zOYQmQFlhTlYFrkCbreM4RjWtfiJEYAZMp1EmZCUbaBYi0/ZxKVXFtO3/
HzrWu+JxXaZIyxlwzQRSsTqcoQSLvCRoYbLKEaAhKdv2QMvLb1/StUOg0W/YoZlf
9S7TKG8Z6GwA2HJ6Wjyt2lhiKNS2LaUSmchz+9AboKyc7GPKGiLBWgi31ekKCZsX
dCklAHvh+fY9HzIfathCCxBLPYBu9a+vK2vXCKOJ8LggUpqsE3ijZ1H9EV/YH5Bn
15htfd7ZbkNp9R62v0KJv8Z2CIH69r2jXYAgL6uWr+41y/X5ceNJydG9W94Y/d7f
WFmTgDMINpskKsQ8UW0hAtq95k7GmBvfsDT1DUsOSMr/6uJYjHIPeooVAEioouYF
m8bcAkYr/UsnpSZJxSqukr1qfGLCz3q5p7hYz0kpe+3Xju7yE04nV8B9jWx/010J
CXY/Z2Il4yR/jYNuGN2mXsM9uSEUBDzOyEISvwYybJHY/yakJUYfX7vThV0/7TNz
Y2xY0iHkzz36ltyUL88U0b3vQQyrcTeHDfnyytw6uIIb3KJI5sYj0DwhnHTQ62W5
inwfcg9OwWp/rMo3LfovQ6nOTmASoCsvmeKG5oNAt6P3BDIxsdm2ewY4xULLB31M
qaufjZnY3QO+1XWBMmQUS2Ivyme9ZbH3NCpnyw2DPVmJ0wtIgUZ8EFpB4TD0lamE
K949WCgFIZGvpztuxSv6HZm21IOfZQxCLN9UwpLbN7Em8zB+BKUBBtgJvTP2SkYT
wKSIqhm4Lmaaf7WvCNxX8xhbxy/kXV/fDLCSYMzMeorC8tIwq52baCpe4VlyUzsF
PHYnJ+nRm3oI2/onSp8LyusPLRah6StSWgFxI5bdCgKARVxuqKajUo9l0TQe91wZ
Cmo5eJnrGNzAsI2h+GWjT/ntfWqWqTukHOIc5oS9SgKNDjw9LuazrTL/n0wlKQgl
feXcdeIBL3mjbJUbzqg8aiRdB30BwFR20/7X4drlB1qzVW7jHBk66RNExuy+9P5B
CbxeT8lJddYYktg4z1kh7Gh8gwvmGS886OcbN+OkDrZa5hWWC1zcQSK/aNgFgnVK
78KY4Mff6nBC14HmqcCAP5JQBPUgfA05lnMzovHX2mNAwJ2ycPLEQ3+40kpAlNgF
RY4qaRB8bbtFtxxweK9KR7bRlxAEq0FkFcdb29jv9EZgvRbfPORDGKcOf7Px4w1I
N9SKiJYn0sjjS3uBYMPUcry+SxtCpcwlhD96tJcU4cO0xBAgQKhiwzT5Trnbfp9z
AHH1/Lc3jIFxtU8f7KTopWOCJ8Olc8a2rLIdrM1Z7803FCpWHRZq5vjGnhEJzKOd
Re8hFREmsHyMSEuD5hnGae+j+T2675IsjB7eus7MSeX6tZds/aUwz14doRZm8+6L
1b6Ev/wRmaFlxvQOP4BiZD3uppMAKxMOZos6GP3BnBqomTetalUygrSbY07tL+is
I1ps96y9W/PfsDha0cdUTX6nhwEyiNOSOENaCAPjlUW0UITSiebE1kye0ZGhd/S8
ei8fbjI6yXJS24r86iUVEgU+5kbP+H8yx095WiFXoNOWmW/HKT8iU7Oy0SIDqLDO
OgoMXgV4NjIIPgI+hcA0GQBTOT6GHlI+NgRmzJ8Li3oiE+JTw/oAiNt+ni1KZ/cF
//H15Cw5YRuB0rTDo104HxitzWIAFHnNVGPsETel8e1K1v6EEr5hVdQpdYTphX0C
LwCV/N2RVS6u164u5GxaBVbJtaw+iTFEYGDpw6scVHS/qFagSo9I0NKaEQda1j6P
0OMJRdEaiI8U/Ou3OKZWb2Mlr8O0f2LNNQV8qbkLr88ht6onnDs8d49q1EF8kvtH
enETrFaWxlnegMEiPQN4/4EJPeCDVOHAHrgkLQm8yHJRPFM3a5PocoSJaeHD3NQA
bSvsGIH0HQha7QKOz8rUqZbkFZdWM20EhVK7t7JKqdwE/D87wolrvV8jtzOT6Tq7
Tm+U0uEQiSAYyQCDTr8Fm1lIjHWNHj37fn46Wlmm/y+CAB1K3wu0PRpVeMVtozCv
bz2pD5OBzK01C010l1gm148e5JhdW455DyaPECeF1AZbJO5DKjRYPpN3jQnlVFT6
YmRcxFGpB2/OcE1nX8Dje4pHdAHrjkzGLdAg2TnF3vfKTUQKIu978XYwI3UCxF/k
hFTVpByUBLNLd3Lz3eO3S9hhnnSfX19VqNSnWysbJCE3izx4Oel2126ZmEgQWV87
x+csK1uyw4QjNk6+ae+LNhFmkggAmiPkD8rTmvcNP7MiC7Alnhi+o/vetT2qhsE3
MAjLT9SS8rbZQ9umayy/Dd18U7A1a2zvVUUPl19hnodRhqN4MPgDa+MCCl9yZmun
4ZU9s+RlvVR9mxhWz35um+dnRy4lvtK4JPvfTEwM8kHY90EWWeSspy2p7+rNS3Dy
si6/zlblvAMLWZ/ijgL7CmWnZb1cSJOWAZOP/+6+48mhl6CjLRgNWmtF/YruytS1
lTes8rPyOmJnxplNm/pNbQAC+jHs3EIdzlpnDYw+MkcOU1KGbR4HRHa0pf481v8k
9YOsiYGkU7focDd0FIEOasqp9lysUw9JlzWnOT0iZjukbvhapVkDVJyMkkzUsptg
mO90Hd9Q57tHGsgBkGNBBmhLYz/c77acdSTQfpd0HgrtpS/ZCIu76v8JyAAKdDQ+
2FbcANiMIpBOKO4liswfbZvj2V0KMgiTAQVx/WcofHfH9GxhIavMfkDtNWSMxWLh
PKjadm4V0v4pHp7lMuQBSZTmVBwTWxnAotERjy5v3Qmvf0L0pWHLrQFPpUfgjID9
HdMmjRucdNLHzMpD0CEEuKMCOEA1/hlOaP/OBE/l0JBeqzXoYRTxouPEa7sBU54J
rXbMl4GEkrVVoCam9eR2Tsqgag7hJO2muW7YNSADxYz1YBGVl72cCAoI1ov2rXCw
TfJNjXcdA5NNGIbpEPJf4mIgHf5Lc+uGYQ0kiJxa8uRzJuTaZokVCW64kGvOP7RP
9n3n8pCaOLRoAUyg+UyXo1A1wwMTULKdpaRS9FLRC1Zj5uDhLk8igc1ZkhDFnTjB
U7Ww6x9VWe0K9riHw1xlfd5sP7PCxzH8I2nylwbXu94dnpGUPZLKskgUKJEKlHvC
YRz5MUZh1JutxIrNfUU6A/oe+PrQPtaunTMTJyQn9UI8U5BlpAcT4l3sfrT6OdW9
FLAftXrwlrW/aWoXbrWDhMbcLNiWmBlHGvpW1lXMdQXQRpiQO7jNFhSn4y8IRoBw
eEXYUmnPuIaHohYhQ8in32tk2ke8OwcluIiMQLpOVos5e94XZDftYLtgCs7W9+4W
Guho0jMyUKGNJGWC69q6+n4XpjVXzbZL6daKpQwcwIr5JXxa/63zCdMZ/quh7ybY
q2zTCYGRGnN+0mxY5IbxRrUotatgwJZq4DUsFDFGf/YwqHyCQbld7tizpXje/yZG
2QGR2wMjwBQUAUwaRvGwZfsYW55yfLsnICiaxhpCIW3xkdoADIM9cRPcacN6Jeit
PuDGLPz3B89z/etVAZB++WMi9TwT2OLiY9Xc5u7cHL0dqrE/mjMEGI+986hvCfT0
Ts+NmkB0i2cIKCpGMMk+TXQR3gLohsiMPnSNmvsLAimG69ehi4WAMKRkFEKazHCW
daRMzRkc44J2OzSXGVrU7XjR+nlWD7kD+ki4/t6eBZeYTHROlVMOv3phUuzbZxHC
lucxeP5Dl7smB57BV6NoBntH8OXZKJOJ7uNStgvNaqEo9491JhNaO/3CFMOKjagV
gJs1+v0E025pnduqv+l2JRxsC0NNPWdRa0Lth20k+pBA35RkT7RNzakqaNtjlVYn
OCv/i+XaSPv6sD/pEImh/lmKzej8mGcYkfS+Zpbr/tbF8yAOozTezfXUp/7igbRT
ac7u3bsa1NUMJfp1WAfqQTScnkN6nVYI+Vf/oZbOhihfOgD4P0nsY8fpkKIhWihF
ErflYN7SYMOY2UAvaZiZAdzmaqbCdCYBVCAhWgTd/T9zS+xEglMI9jYnbMGo7o4z
AiPbyAmQv5m0AONpAKV+w5g55Y1DP/oHpFxKZuJnHSMzPKSztlj9y/i/HCxbp2p+
ntwwHU1iJfoOzyP8Nxus09OvNcEOO5hiMRABI32XM36ClIWTkopYq2VF1AwAOvmp
aU8tOBD9+2G4siu93wG/RsKcAW+kaq7LRYtRSY1V1dfY3h3rmVPDq/FtqE0gZ0EB
WZXtaz7S9SocvZmtooCuVjNcA1f6uZCO0H6jvICbzRp2wxut6Fi3yfeywOwRQph0
HpPfSkUN4sfCpuK9LNLoRliBPev3NB4A0HJVV085f61MD2YgF8o05vEAeHbXn4Dy
2er9QXCj0TeQHs5cJOxmXgCbAux1aNebcHd9mttp4zdZNqMveyi3TarFbhr9dXb+
5zUf1jnrm/QaZhbjWCb/BD/fh39ZuQCSoITwQCp9xZv0Y8ab0Iv7KKEq2gyfIGZ7
XipPu1I1A4tvjzUTuRDKXiBeGaX+6aZyj9dhzaJLn4hHfcrMptN61y3+bXsVd6ad
8O8lN1FOfurHga4Yi89DowbPIaDIRx4fRcqKqIOEhe1C68Petcbt5+CzrW513xVi
FHuo9jGprgAKKvp/zZzy3/O3WZ6BK/RKv6hMsmO6SifV4FfMJdwnztvs20sdmZe1
nzhXDIZ07wg4Q/i38VOCBtIaGWKU+M8voMpoSkEqmhA5+fYtETJIlkC4YwI8zrI8
/OdFkstPnmxddn3g+SJf3BTa3NjuPpelJaD4ku9cOSDoGrvJd8QpDi++xVP7pHDi
m1NDd7gYvQ+twSFFOkx3iqmu6EO4lliCCegEQA/j14AqjXMTGA8gOOCFu2ddckTE
6GAhAhH131yxGIQN1VrqVHWsz9emLIP6VHd4g5Pe6bHjyMUJRSQzaqkgttEJ2ZoB
S/KzlqfRP2yo4LQRLVEfVuyZSdiTzzz8lv+rJJ5JOq2IgJxXtjyDCkL1gMGS+9+x
UJOe06uUV6HXQro0ZRWM22SfHWZdUkhn61M2l2g7wpUckIqPptvDoBTAqHYraEQB
6j72zD1LAvqIswLQ0nv1IXqahmExPmfAcRpdtJWO8BcMMAlfJBs+yXxsQcFkk32y
lu0QYWvK+ZIr/Rg8rgY72NsoSRPCK1g9Tk3ir26tuUPXctE1umPQXONKoVfVXl2/
eJD2SkjwaX+eJv66c0NF/x0r+3dz4xeR+7ZyEtDGTlHOLMeHsHrkMzi7wJIsAXB8
avkOJDdyYMtYzGBAxGji71FbCK8Xh+/RxyHAWUfQwtpxKUXIvBjqQxUXfprSinNe
zKx0n5Q68aymrQM5A8fwY08xFgu9x6NeFXYl/O9p1IVI7unq3YaD7IWIGNBzkra6
55rsfYEJrPh4gDNLIJggVHjoj1AIukOEaG4P/mauJomqofOUZByHa2N/BDS5dvGL
KKyV8DJ3ZXWiSkVdp8CLMoN/7M1lTug2Tz2e6Zoffde4ROUJgr2HeBhJainx5mJG
iexTJch/WwqRYsQwt99UhCBJbWOJlI4Rv1xVy/XN8L2SWdoTIFWcQAjPuRisvAoG
4orhmt9QCzgsus6QnsbhXiUoJQ5HuFi+krnazu3eGHAMDlfA8Oma2RcuhtqCxo0t
ti/UMZu9LkzzX8z2XIGbKrabMVbkIX1JM6owehVWieaX3+Dt+n731PbWdsZMAzmO
n9B2fPEHacWn6R+wao0IvfjW3Zr1RIFfQXbZ8h9I5mEXc4COv2bPG+mc4sFTVi2q
spMWV7038UdEPSKuEHEULDo/Fcj+PzB5uDfRPSYFQuVRqSyplXB8reRMtFkZPHZ1
PlfTUZKQlW4q7sWmCdoeaImrtkHd2B+80YS1SfhYljF/dq9ujnVy1z53ZomP+xF9
+bikOItBVaVV3QNXRFZVhZkhB7Z9hu2iwt5p1AC9QjtD2590d6NrNVSr8Dz+OE3m
gFh5N5bxMbYb1CNZ3plB3tfJKOtceEGHhPQM79zvgZuz9Oi9Z5Na741qDlw5UP3B
F7RinU7BalPmxCrzq0e2qVXI15pdr4BaBFGhsQsBtopRykmGEoQl06oF9cCSO0Ep
DWvxFrRsKm5afgUr6sClkCrjU2BcWAgcInKXoQaUzajlh6+5lixdB+7bJ4L5UElQ
MHpgAs3Sfkf5dhe9kZvIq61ukNEcxzaed/V+vHpMModzm7iTM0ZWpALD+EB2xB//
ce8SFuXi5/UfyAjFKGTb5H766kksjKydRbWD6SAhcI/mX24FBr5z7BFy4/Mr4Va/
rHB+mcktRmH2jYunIoj46W7aMxhNvekm8NtYB3YxEZHYT6NSMeu915z7ZmaJv7Fo
KpxagTx7GKXcdXnF5xRiId5ulHzK/O0Vso7CwsOyUHpqyyl6nVY7pZN1H+J18JD6
27RH6cFKWS8GZZ4BvHnFFn+3CW/P9R40MdOlej2x8ZyDnMo+wOoIe6jj902Z4mhi
eRp1TAMCQu9Hw4KnFHEVctJCXUPdvY2hijZ3p8DJ1q1K7YXkuJSSENWkgk+CHE+A
gl1DigLeD6zwh1926J7GRCALLBZ7k63ZpppjFZxLT2azKw1VMtBnTuW18/0sdo+A
p4z6MpKM5lmowecuadqjCZ0ltgfL34uv07Y6tGCyF+TAHwtkw/7/zi4zJldn2pfF
CEpK0HPBFin/apqQ7V9UDk1jpZuaAXdvFq7l3DMyhZlMrXxXCK8FTMdDnhzdbrsq
xMLhl9ZA8IHcuB77QT/mDFkYJSzia9HICm8akRyBIfHVv2CtPMfSu9sYbuRN1gEz
SdwinDa05+mTuU2w0ukTY8xSs7sa/360dY+yFQ4tn90N+PaWm7v8VG9Kped0Z9DA
QesKXbTnQdhv9yuxJnuDs3vlgP70URWc2sLEmJe/2L8YbpvFk4QSEQ7DsA4ZF/y5
qQIlHjeunRYPiKZXKrZPh0apat2UzT4px/v4arwLT7Py9ST1CVCfzttXh+n5x7EQ
3LwhF0T5bO9vaxPCYBP++LTqD/qGGeRvG8CJfaftLDBTfUbytgWLNkEZjyh7UIeu
CKJJIX5Mt//Ax1jBIlrdvOLjxVd760urFDoff5lDDnFVm6k3zz1vR4GYGzq8mrRG
0g4pMmBB5Ah1hmsl7NI/vYIJ20KfYqMaaQbmk84OkHDtlteaPzvjtmcgMGKN8WKb
KL7ORhnN1FE3xJ9fSLlLbIdEt5QY8v0mp76lRyMXCZ5P2JqRzXJtONagid9iMZD9
R8ioM29fDjQOM1LVjQ1a1GnR13+hMnNZv3BQjzqPjc1tue38AGdgR80B1p9ztgfs
5R6ZMjLXvx6uUDR1C4HQJRpKZ3OQddjH2eA9PfQUveB4F3ihvS+JW+H4oDwpukZ6
OJW4lNY78IiwBe05r/5vz3gDogudQiASxggZY6a9/RZ3pwYthFP/BP3BQ6EMZ+zA
1pJsmGRgE+zesLk3SJQzIVSL9XMEZDqG+58XVqipSIHt/5AIscpqzNxilgMFUbxp
oG0+RiPmzn7FdzYFEG+EEZ+1Jpn4fC2fSBY9rCOxSVBKfUgBn6Aa9luNOf/OdIUz
5hCZvz4PFFOiDu/WEGSULx2DlCrmWkXPK7/DlEEX0RV6YZ6LiUFfGyKYN9MUY17O
DMrO+IM2j61C3f4ZKq2JImsLLQn5oe24lDBnd8bT/ojoEin6s2nZW89e2BsPh/yV
e//HKr3q17HgfSLTfOkmmB/BmvXXmF+AZop59k1HyQVjaUudvGRcKBtYeNxbWfcp
pbESlF/oH7S7+wxb0CfHXWim8931tG2eM/XgUIYbeRcemT9uVp9cOtnOCkJfRaVx
lGANEE+fYi5ZY7tu25IGtJ+kwJNBslGEc0ggc77SNfRApUN63z/mibutNK+Bye9r
sE3y+oASITwfLTgqiilnb3SwW75xGJPx1gEK+aPCMDqtqqmgmFzGn810e9XEITH9
uQ4VG/Sf2DRwKnDoGdo3JtbghZyqPUF/phC/Xq2+Fg/kzn3AfrVNXzzAYtyuc6a3
xh/FLZ+TQHAhEvO45tUOIJVc7wklBztgYKFkTpphc6t8pnFySPdBoDmGw15DtEU+
RsSlOFnmCjBzMhKYII8G2+rj7wTMt2GNnK6yyGS0ipwwKWAzg+aTl4o4pc/fYP/M
BQWM6x4wU7Ods6PCi8e24oCI2cFEozP1qiA17MK3SZKGr0jX7EdEo02h1mbnMkl/
cuqwdTg9wzePhDYPomlKV32o3axQYC8jNydkvDWYU22DRQtA6mGNqQwIXsoTPkv+
XIskKgjaW3zFJ3O666i7ZiQHvtIV5H/zYLT9gY5T6GmF+dsg91TO92FKLuZBd6tX
aJqHvbetpNCNRcGJNIDcQEHOwiZ2NvYmSBfXkqLHCPWlX+67zkx2gHiMmLZ4USzU
u5PYpCG7DLNLbeg3hNzZYBvApRaQFQIz5cj8g95pR89090qwuWPqTB3v+gMd3ry2
PpNfvtkVcibeBz099RjSomtRcG/MzZAcnVr+emUtwwWVZgY1DkFYZBEuXC6NXfqn
/d+FQV5SqEYL00uqK4+BJsXl2CTCU8H75THl815FEiXBm3s8hruGYWE9AHAoFcxA
srCmcKovEUtW/WMlwjkrjOXv24pT5JcnfOe3aIH5HwnXSEdCNbxYYGQkC8ME3OSY
3sGfb5gGtcej7s4XSGSR233kt44tpwwuC9OVcsUfYOTlphjyqr74QFadL+wCK8bD
+lFURFoshCCkmJ7Gc2Z2gWMoSGSx0B4W+mw9KHDsVJXMr2D4ja8UGd9+Axn5IAP9
S4ugO5UgmgAIvfZUDnHBcMZOPLDUzaCpZEpK7euXXZe9idKWXxHB1209pxq+Dlb5
dQoIQ/r47sSRcyydH+bGjTgT4hG2gHD+jsvuG+4Rjcy9d5mst4p1T7S8H+ZWmlCi
0wCsj8h2TqdTSvopE2Eu6ZNULLtAVoBNoPY79ILtPsQ7gvEjak2/lLTfsApHrr0+
/LvqzlS3tWCQKMsxy27iYLLwaeLbFbyeR2UwXfxfdUULP/WGtjsaYZtk9vxHVS0n
pXqRvzrqTqqxfQZFnX/VjquiAznJYJPkgsUa1QzWifSGX1VtQvp7dHTXvJ46IUbV
C1qM8zsbKJpz7UrBqiOH6CGJHSqV8+AU/WrMj9yInZNzWCobHevuRW1X9MHfF3zL
GrHr8qX+ceOSk+6RyWFfn0g6gf2kel9BKP1cj3oCurZCsGEHsKqJGTQURRWYo71E
JE6pRl4/1fRJypFV3m+pd0gZXVhyiBUWlFEq+k/sMWvaqJnHPbJe66KplyfpiTZo
noJ1WDKiHFCFuPmQ+ttqT0x9Yu4K5467oEj9idgzzh/jx8u8cTzzpB02SQG1avr4
UwmNO6+wkr38BtztR6pFeojFSqgEB63lVl0ftgMcG4d2UghaEX3+WOxVKAMHrEsn
mTzkT7yPVVUfDFr9n74PWADrQM6KGWdDAQqhgq/Wzw9dYZlAP96bUKcRMiZMnp76
F9BWRo3pWsGlxM3rVLcocR7pKQ9x5v8JdmK5q8ZIO6uDobHcDfpyKSgVqwi+CXeS
XSYLT+kpAtasLnv1QdO5H+JtqrPEoIE4uiLYYjUEsRacZSiIWcW84wa9I6y2V2VR
tMcy+sDui5c02KnulCtArzxR0904A2D6xG4mue5EmbS/nbYH+UF2Fkc48ChKL87n
xVUBgzDxk3t80Jkj5liqPrg9+/CQGp8ZFnct7AmL0E+aq5+OH35D6ETx4E5/nZln
E3z4moNv6MUr7m74vlre2qQeVv/6RWs9WJnbEOJM92R/Vp3PI3X5XO8gBQIMFFYX
3T+qKNTPiRzARALhelM386ude8PbD6YFdsUC/txlYcOK9sZtljWb6JI211/DepZq
Fibk4j026HU7TYo3z6HhehCIG6qW1Fa14/oRgGcURwJLLMSNt0ML2ZAOqqZx1aEs
NNqZ78qGK/ZuFo0mpb/w093XENPi5Xb9WEcGBdT6jxp6kYRUJ8J+LqBV39o1kHUf
4dXWHa5scvXvzz9UUqJSPSfKUbh7gwqfmo+UX5q7uFwoQuknQxJgoSmUGvByTSDm
Lu3G6SifAerr4Ev5svZC2LrCsQfT/P1Ee0evaL//es+oekS+KUSlgnXkNRSMTG7n
mII+Tl1cvxkXRBQ3lP6vfkrMkAy46rHFAqqGrIYtnM6uw9vJ+9UFRrO/4z8jG9Ey
0OSyGYEutJ/wU7IlyfeDJd9PNTrdIKTwCSXwWdnJ9J6jsYUcahYD/Bv1npG1JvGU
cfNMEdScaPIso76ZlkuH9HBGzf6HCf+DqQ90Woo/Y64uuY09gh1esOzQGoozUgrC
gKz2U3twWOersD06+yZceol4eR3fa4ZP6o1b36zjxmJBTpPJ4cI74IiSNX405Pm0
6DUguZG7YmWEGhcNN8LVppLlf4TTYLk5S8Z26cF4imlqbcLx+9RhTOJM016dyz9O
vp4OUgL7uoiP1pxqk7cwWzPDMPiG/snUg0uS7xc+E/cKhwrxPSZdRzJQo+q9swKP
pCEqG7nwPZn+wmKaK17qx3zGgD5NiEQ2TaOUvbpp7fuEx9Ky2EwA3t6Vjw6URlyM
Nwcg1h86l12qyFI8JatG/PjR28q7S5MHli9x4v9aVcrgfIh/BOz4ww/R30TNbQhU
AN+7t/wYrYg5949l7/PRra0ijYbYUzPqktnyp+I/YWFK4aM5bNHWQXaoFBgXyZZT
5RooexQol3JV7+dtWZwzTdQark4UWWg1dSwXTu24B2EL9OEZVIi3p6WgMamOL9EO
tSk/KbM1Npc00YG5amr7itHNdHWAkSqZ3Fb9nj7E5zFN9DM1lOJPBMAOTa6sHNbP
WzAcoU0EWKYVQXbY6YBb82Op+tWoCMl+Tp9XoalsT3eCQF9wtjIzy6ChBl50o5JQ
KfkzcRSvvZpdsxrc2XjASVOh5NrahOSoaDKAgtujaPfC5KQX/zS30njrhKsO08F8
m4VSzlZcQOtM7qiG31xATV/csfWWkya73y9djd5ByrIw1REJNzuRH53pHbaqMEIf
K2Zi1/IxVGUgtph8nHQ1ldF3NNvfDh24Mn/gki/56hxkWKv/SGr4zIGMIXpQLPLg
wmSg7lECoC/2L79lBStPgEcssLNK5aXYtPlYcIQLF+tyxiNnr5LuosnQhzvcaCEh
QPVJtL+rvbP6ccvIzm9gk4gk6H/dB8LE32YQeKN9Yr/D8Sy5TTm+dXKMrv9AFkXw
6B2P4pen6KlbII/aQO4frofBUU80dYflWHYdSeBtoC+wOu0ZYhquNdRqjOo/iBX2
e94jQMs7wF21kmTIFf7gFJjSY3Z1yonqNHmzxNqsAPJ00Nah8463WAKj6oRrfej2
DLglRTlQyYtpncGhxgGIRa9pL6t9OeHKD5cihz0qpyxhGl7jxCH1VOyeEL0J7OaX
x8QjMsiJHqwimCmv6qYMiILtx8uLj1s0AECEojmDo5CiC3KdnVrL5FnK3cifdWLl
voXjAeA1d8cAopryr2lPyef7w4rJbkrpnhFhr4+hHy4yg2nLmyzok/P05Wjs+9IF
rxNcDZGsgLbsyxoRbumUzoEOx1TA27E4hB0FBTNKotdi5WLZWEPHGlJDLDiJllaG
oNhRrWPIrGgkYnmE+HAlurX3oNZb04dniOvzS3X887TnSXO6p0qYu+xdGJ1Z8jwX
Z71ywJoOI4G3vrtu6W8pHiv7gtMJANRgn8kjZM+/JpplNQQyt7feYmdx5wMknwPP
MaE6NpHwdExtqgnHnBqQAeDQH66CsX8fFvtDI5kbWMFc2ctxmCOBZTvH15jVip3Y
6eW8rRL+8fPmN7XCEAAsAK9TFWiv+VsWANetgYAmO7DxJpsMzVybxe76AjqapdzS
cT4TdTLfSF5+TDwm91RuU/+nKQGp4m9PCr2kvOxvx4cuCMCme5bxKiExCuZO44WU
Sg88M63L1E/LlnqJn11MUDMmkdjbhk1XLnBzg9EhB/dDL0GWJxNscnA4JiGY4UbM
Xd3UYxlMS2V5vm4NNd/1UqUmRiiQvjtLnVw5j6jzHPsrFJZHTig3ArQZ4s7uir2n
TKz93Uzw2ieHxgzsdqsolNqbehY9t7QWKBgU82gt4dslX8Ftv6+z1YOzaKbfMjU4
g+X+e2P5DpzXSNbruZh0a28iTCvA5aV4voAjM5uVR9xl0ZtE82fKOPzdEOdfjq2A
JF5+LdCJNfUGaFRCtDuwYwqvOoHIzgBc8mA7nOnoi9Is3KUmDXYJtkPU1EmLjlVj
jMqrxPFBcM+vamB+IHx1ItUt6cztj4Rd5N13eCfVacaBzNa7JounUFmNuiK49Ox3
UnVt25HRVS2Vr3J9a25fmzzRv5FlbwSjHjoPLrfMPjJgp33LKrouDRNZNLf4hCrk
R4vDBJQNAAeAiNL2USE1FalIyCoN3H/q/Voekxpa8eBuiDtWIG8MLp2XtMjBzbtb
K8bPi9SUMhLtA0h2pIDZpOCkK7H8B5VQAdRYsvvwCn1Ig/PQunRsHMciej/YTTSo
SuKYEsnNkUiMJZ0Em6LfwdvZPTVkfl/a4tTO2fweBuzyACPIe9XZ+2Hg16hezpdd
n/Xc+dAG+AUULEXMdjqO8TfuFBUhy/VqVeYrASicjFhttZODav+ohplQHlUiEfXp
woL8mVyGhJ9cXVpsYarzCS9QHB9Ymy1/f174wnQWik6+xSIdD+HeFFG7apYM9UiE
8QYWUo9sRbuToyXX3aYAQBCUS4Fr7Y6/mU2CfL3BcYnoy96NSB0CCjyluzH+xOYW
FkgjsEaNdq+Bh5WXIFKlCBdO/H36USqdBoJqxnMgiYh8LTX/yU8EPic0R6/7y9OV
4oTsJToDQKs+izXdwMZ/wMjmroGcEAEjKC9ObtweCloU598djO5FBdSvsRxh8lL8
fqXUJyrDmBWuKDkRS+nHtCap/rAiPUF8HBZao0au7DAT0Dm+BOl9QHAEy/5WKeT9
hWGy5yeu9zWNTymq5oQlOPkrp81Hhc9S9c9yBDukA3T8dyEg7cpkEfnDF6AQrYX6
b/OryQguBXaqYElyewtbwBcOu2yuUrmU8mCZ1IfyDb1AQyjFO2eJD0X9Krgz7si0
RD3/ed+Az2lKmxwv6DfQL6XZXbz0BpsSmG7WI3M66mEcI8FEJTdlvMwd8/CnBt3T
jalF7fuukr+Zug8S4YYIuvXkZ/wQmBsW3o+PWEyD/wpTkimBh8ZDGsyGi0M8tmV1
oIE94X8/umNdQuTu+GMigO4+Tlh9XMKZ8d3CZ9BOwhaP1a+Lb6FGVbDwuo5mcqSC
WyOEj2cRL3VWzGtus1IjcUaOENCaKTf+0DiEX7EbcansZ36PX5+VV9m4GAo9I52r
6k5WElZDpPxLD1/cs/DhI+qGDOpR4WFBoy1HsyRoP4rWwX2uUH4oLwjiYZ0e3Q3u
OJxovDgQ7Io73Oc02crakdrkrTKRYoQVsiBSuYxNfN5OyHqi/rDhuS5USooCRKOZ
Yu1IFPrjjhctOqKfQL+PumL7zmQkGVPGaza7dk7R6l9lPMIbHV1PpzdyKHkX3blq
JqYpb1we3Hm+cefgzSD117crUDgbEHQkru3x4ufEkCcBnQP17vL8ja0t2t9/xjI7
hwVQMExRQjiBhFQYnPgiR5P7i0dsCidhygBGbAIpGKJY/QD+NOl1ajvmlRWtrkO2
Q6oasxLRh3jmjAXWnr1M0vtVdI2Z+Rq0Y011MFykhwEsVye7ONICt4NvJj0Q1wfE
HvMsYHso9BotyoEEaOkYUiw35SHzo+Gfq5EKEAv03dggVx7I/kgeWFW+dWlQ87Cq
f0FCREoPL2cXvdr5LNcm9zey/SQKjza5z6v+0xKpbnZ314jeuSKMlRSJ78FsEFnj
vjRMhn50y1hQFaKxUZQHFVWDO/gsyi5IeumhqkyLbcahTvIYWHBMgMP1k2Aztgfz
9Sy9gcDOhmvl4PIiekEafBQ0WQ16hx9n9E96gSIApxKjwfanmyVSW6s6btO3cyeQ
mMmf6egKXIzZvo5iRj7bsCXMxPWys+vX+f7lA2YowcPrpjGGREKEaUOvegz4xGgn
XitunlAxdbWJCLfLNOJHQ3Lk1D0MKA6kAQGqJKTBsNOK4W9H2IX5cUMjNhwAtx8U
JNlxoyqzCENrtePxVmE1MprPjzXGeyh8iBaJy14elenlzyJywqAk5cE8+amsgBqx
xRHpAaHLtVShFBW8+oNvzIqj8N8nF3c0yrefTD2FIwDQXeZ2sqDZRpPUcT6SGRbb
jHZUUoaV2hAxLwggcAc30Ab4ge+CWdEsKOkPmk7Jq3GrcHPFPsQj+qhGdWISffUr
j+zLuqMAMAJvlNvEnC+tPUPiOOnDj80urBX9Ypgm65ZVejIAOZhpq8qprjup5F9Y
I+THDfKSyvJWn+RKzKAF/NfsC/vcUqDcbuR9QQyTHFiTzbIiyQggUsO7vziq2rwA
A3I/6hPbAEdq9LVQDg67Sc7D1dgzGcAtsRdTvMQHeuo/WBjV2arZSsCBZRjI4TIF
VI23ufLzwU8TqMgELTqT+T4T5wBegMOBrJmbzuZ/whLxxQmxBNMD/ySAlucnP7EO
OOLeA0sbpVX1KrUiy3L/3Yz1nttB352dARlam9yQTkkdETPssDxktC5bKopRpFI9
pL9SLtJA3TgBkPQ3NnxUH43CfPZ6wpDwGsxz4DTISAwzUM4Z1hgRqsKC+/v0wEi7
KvMBXczxU5/fpqqfl38uIX6lY91eUJ0o3elt5Dxm7U75iIimiUH64YlDLh+tkkp4
HhpQLMawtjzbDCyWfP1tfzA3N/1Vq5A2+PtS0wPpUqSS2r4DDjrg/tv0mKsuRcJS
7doorWBgLiQLoEsfiu7LHwUapxAVTJg62XZECrug0h4nm5KZRTLqpD/94fiJhJE4
giOvdVFwmBSFfpGmhEl9G6f798XQc6D+rBBTDnZtYbj+wTvJXpBKQ2SIcRqyTI7K
RJqD8GTtdqdYdZZ1Ut+OSwRqx4erkIViyKSo4YKs+aHFFmh4a9MQCjbQQanvoCiS
R76K2wbwCHjXZRHJaTQqPDPLZBssWpt5KeYK3cicmTWDUMJPNcri64iNMC+XM36r
sQYXqBa+MiMODDbNS6a420gIvFH6dFbAw4zUpANrO/Mgfl7OjJ0rkNIxUacF9I9k
5cUX05EsQL6rhj/zOfC5FO8koifhkb+ObzWOK4HncpepGgwzmC39VR8fM+8WDnLa
REr5nkK1kJipiebZVHfQQD19rcEkGuk0hjaG4u7T9xrCPBrpE58U4W/Ca7D0W93E
E+kKmRwpFV7PaGdhCFhTnVppo3P4iWtGnxYuTL+2F3pyepx+CmAm8C5ZAe+n/Nx0
Hm9hFQWqOgInME96aC2FpnX2CkYemron10JxN6n6hsB0ZzgXf8auKa03V2K54kGz
vHSMVqNOfQHfgf2uQx2616vgmnEXZPaPu8mvDYxuxYtvFAJz5lElEntsd7MxaY4S
Fg8twx8gt5bA0kokrOxVCrGiBAYu2SpW4V2ZOUj5QHW+MXNqqARqFI9eKc+p3iCG
objpz4geRK2zmE6goJtBtQdq8J1dgKyYyZdp8uwG3lhh3ozPb6EsjMxM0DPRuMf8
oTeu15R4FfHALkD8lFBgMKShw7VvlmTuFztiTsSnwJft6nBX/1K54kSOFVo0biIh
/POYlXrDBCMfeYb2iuvcfpZL400pKLx7J/hlQ85rXTPOCO6lSL1Ogt/HOpL9TZ98
i2lQ7fSyza+K6DpcHHB0YNitN5+/+McX5vX0piMiC4S0jBo7y1QgBfNTYd2TJM9F
M1b4d++v3hjXJg7SvorJqCXqwnvrDRRqKqfpX0NcmI1JSvrzcOc3IRYLLKf/x/ZD
/6byyRG13LVkOIsVRcEjnT1DD+3X9KlD/Nuo9u4lsUYw/P1HB2vQXjgxvDT9VhBm
2/P0xHy7kMUtdIyBmZ3Dzg6bbGDUZ9VEB+W6d7KfeDmS0IU5DItk4blYbNuZBuzr
vfWAhcUrqg0CLuxGGhGi2imkl6Y5sDO1o3S+IFOVCePqxFr1Vx7YNXXj/9/igZYv
MqIyt38R90uvPh57qI7zeOaocmno7wQsB3wcVv/HZ96Sg2ybneCrj0+hdFHTzaG6
T5Rlpblm16kvSA+K8r5OtDcHtOCZ7+8T1njXPajtRqBk715YZDLr4eBWrGOVm7q1
9eqtEAf9KbBLVp0CtZDq+jowZAeJyZYmYzWfA8m7JqjDgRz5qxf8BvIV14poCw6N
kdljZydHB8oNh4KPqPuC/iCdo8vAkqtGWgcn8FYN2orEjVX2ZAFxlOJockUB8P+o
8AKBQPn9IjlhT3eD1l+oe6AkMHoqAEG4Yew3qkJqBsmp/vkNwBJ5PYHa1dezME47
bNF8ZcTBZgpDI9M2YFQA4qT2FO0m60pJ4Gf3krqJdMpId2H/4n+0iO45afmMuR++
pcHithmaL0Rr1QGtaVmN3IWyzWrjAIv2eq6E3p7bWN1XqNRfKPDNBl9pFWmkVk9z
k2FliD3NG0Jqn7mxpVNJ/cQvrayz3Rm7GCCG+rU+El6/Jz+CwKUr+ImWfNWE1I+u
hp1kkt8EwvysDjc2A2aaWWhGmpIgKeqBEItkCBPI202AH2sxJ/7Q4HXr1Tx7xmBo
6BTppMG2LSvD7I/BMtEs/wrgozqSPkKMB8k+1+Dt2lwFgtWJtKc/L878qwEl6R3e
UgkytOZoFKpBpu8vnpLFhJrXnq+aiXoxJ4XDY5wpQ9e8I4rC2Tq6AEg04jyD91at
9ysZabt/cHHX7e5hiIzJtco+jUqQCcIZE4WDR4/Wl2c2HxqaMeIw8FguhGNE3kMx
xYJyFBdpMWTvWaSmF9pj0JEVffI/Qamoz+xUC1/ui/vyTSZ8kTLfla/VloiW+O+V
vZb9/Kizx/8WG+KNPqXG+H6D5GjZAJ8dWC2xIIjiGfCBCw36WM9t+dhq+iO6vd1f
2tTO6Zb0WoigYy90awbFugoQGMaLkw3cQCzHz8BSee4VTMFfhbkB87CFDHRkp3q2
43IuQh5wG4FVGlGX9s0jOTRd7J1rvGr96wuPXYXhniEEAftS/vVO3wV922O0U/Kr
jt0jJisKxcWSzOa4vWvSJsdUxKdAU2y6jybLnEm4l7/RSLZ4VlztNe1JJTpRPiZy
hwEtusDgX5SPn9SU4R8TilRRMR1obRbSYwOh4qKBBPVe5SqpllcHou8iDu3sSeu6
vxamF1DciHHvbZ2+aLlRLu4UYwnPHMo5pZusYRCDQZJbdBYiXW8mahKA9Di5caI5
fLNVhVqqrz8I2lk0MaqWA5mjdnKp/mG1j6n28KWU2SnEI2+ZLHZL3GqGJPdRxjPB
FFTm6//DUtdHzNuYQDIYADuOkF7HjYv7ikUsffdFuOX9YTi1+L5731LGE1aK9GgK
CvIiVMz42htPlU3nS/LKlAT9wJGqD6FZ4mEi5DORtK6EHJZrmr8aDVmr7N0a/9aG
dvaOY9ur0in6OIDwzFHep2FwvCmpnWsk4iRnSqdY6Twqmb7KJk5bNVAnEYuCIgir
Ae/0fOzwRRIsvT1C/NsZFyDBwgi9KY6Mu1roZR9wbqL9AUdIe2UI+bF78BGXSVly
r7GozJjLcDuMl5GFU+rYaF1hEqwdw4LN8CYg5rapcyY1R++OrQVnR28V/FPzVY1V
KtSYH9jD+4dEc6P+Noos6NzWJzd2Hu2HTqloPyydsThwnY5PlgTg2wdWP1l8DZX9
IsegOptKEb04PpFKlKK8VOU0ZnpCIxltEsdQE8OS5R+GbGj2oJ6LODqm5YLRM5Mq
d4C4zD1M//6gL16eXG+woXAD7U4YwwhuupB1vAZWwrJDoUaMQYbh82sLrmTAhGZ8
URE9JQf56h3zSojcBzoW0D9dBged+fEIN6zpJFXCWMmyoIijpBiDB3xdIzKhmEwj
0JiMoDOR3swuhvv4PsN8mdwcLUr8PHsLvyu8TQAE8SgdV8/dy3En2VJz7TYA8leL
A2j0aXHfA3F8nHoF5EueehYdzSfw9GZX/6r16JmbH4aMfQT4fMAd72vo7yFEcYq2
AB7J0+SmdoyYBHqHYrghrYy7oZ1WP2fJQFzqqBhAuQl71bvZ+Q7anREliYjAM8V+
lHRwuVpE6KvZ5nS742aCVt8yeNt6WkpRHabCuwUXdvK5npsjF2irSTyKXgJ7wo1r
aTMV+rdEGi9b4Uk/CuwK/P/MhqpD3Vhvj3zOlw44ikjMm7cGta/XbD40vJs0ZSzr
oehZdLUiYAm0bhJzGgjYSSwmSLJEdOD8k5DX+ikcC4yvCPRDKlFqE9Otq8PW8bnp
hndnA0T5XOFg8DiAZTFYPiuAinIjbv70SYr8kquhSBfEoFW6SW1YYZ2eQDpzAR8p
DD29zXlIuaswwpzjNOJaETSNaY3fJu2ksOSNHSeqel0gEaqS9anvnC4OLK5RumXo
lbEbA3vksyzUv1Nh4j6h0avYcZgOEJDDJsE4Zejt2V99I5d8KBmBY7Ic7hLvsL5A
VW/infkT90whu/aoItIOoYgCerogtyBpwiv7vZis4HfJneKC7Ng+T7+M7NgsP9vu
fKoSLK2T0F80aVihmNQ0F+iR5naHq9g6lUVI8VxMiq3bBrMjDMK2ytQYUShtBX3+
ddsV3O0A4lSSPeSgM/4Nv+3iF5tHzwg22OAgTpc/y4iFUziiGEJ6vPgyTQflI8eE
tkfm2gA7CqmcgLEf6AQaHApn1q02qKBSm3CT4hXzgac25WWhFsMHPc5Ubvz913aq
jhy9a4ZpvLkRz6Na027svZOkrvuhpIibqzj+MmE+XvPrVxos507xWWTNYZv2Dy27
grte14cdh8lXblnhsyVcAtemgKs7fCYoClkHNaBNKyk=
`pragma protect end_protected
