// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k4XAaqyYhBebpBHzjbJcGhWiDerckWdKC5VTI8XJpJFT0ACz1OOLuGiIvGoFNJIx
P4Zej5jCpmR69qxGvhSbviD/3V85/xGP0Fxme5PcHPB9ody7kNfRLwwZFkd1Yobo
c46uuucqTQHAcoGGdV8Jb+80VSuMgxWl65mSRBm54N0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22128)
6S/KtKJt1m8kpaMPEhwyMNr8hI9Eul9wIlgsqVqbXCkhLi0aC/m8WgY2u/TbLy7a
6NAhmFAg8P47rWiBnWZJOnSWFfo8RO8KjTSnOpveOqg3tff1QDQjdeKted+S6RBP
Rul9L6JrmwtmgTjHBLRoZ62B2+GevWCkVLQfMuuAoO3ExpimCrGEyPYGteuH/ToF
NllcjX6wmFaLTRn7Y91V7dIs0bqvhJ9/E3mdUGbE5H/h/k4cLSKoiIAKyJsj76pK
5TROcx9SvM63wI70eKLlg/6AYhzws7qDMgYhJcFcotFbSCIwuSsftfHd5EdDUKGy
DLln/A1dYFrG8LK8z8tO0iqSdriURDX9aBjIfOLW0KWiWgBPWXppF7f6zjJpHu/1
JthVVvFKuC/OASF53h/7YA8aYfDcGcC18jb4TEXgjgbGs/mKr+VLC0+49+lWXXWi
xPyHhGn0kzm5fv6WxgCrRjV20pXtH8eUB7BDKLl7ruJA0+ex9wvr/Dq/29L/KDEC
EEhTfNTaEoAT5U1UFE1JzR0j6QEpeoPKfCdhChUPNxbuQGLlbkUmgR++z0J2JECi
J71coFW7JOt8vOyhSfIfzJQjb+Uz7ICFtjiRgKIM3Y6SBKofkh0007F5YXy3wEt+
jrGGj6Z8RQO/WWnYxHQRWkT3tPPmTa4OL1MMlPrmu2eGkE+AiV9/hEc0m6a4uKUs
xdUU8eTUCQAd1ANZ2iQ05KCPucCYhQkLbgJmCI3WU22BQ/7+7Tg56F0np7Rch3/x
OgHnphTwMkUWnAHPlaOlD/ED7skB2orW+eZWw931UiOZkOIIA1Qvv6Ebgru3ve/M
h78EOb3Z8+h2hKXYDcVrQ8Sz7BGbT2Za+tNGhM4LXGVBVt3U7kKNO9JQrgNrEqc6
mMQkF0Ou7AjmpbQxAcU5d+EP1hBb8hE5CEtD0ICQEOxUMa3N5mDyE0Pzpwp1Fc2L
aBEMJfke4FQh1dqXoSYZXDHaJIYnrhzELWHgFg6ODF9eB4i3mSfPNke6K8yuugGO
r7xZuraYgAolhLQ8OVbjYOAsCnwAV2XRGliFp+YhfWtchxDflSpd/O7vWNWqxwfl
E1dY1uKw5bn4X4N/xbGsOW6m24SErPV3Z6UUh0UrWxgMxDy9GBrq40RHP3DvaaJj
mGANvEWp182FktLtrLd4on0XGFZke3h7nkN+N7oWSS5vPfydAdE+1Bih5Ew2FaO4
F3r7abGxMCiQTI0YRgkW3jLl5huX+JIOPlQx/oSMQDzchrcrc27BcKb8Pq7YoJq1
V8CbTVWsPNPG0F45WdX0iRf96L7ute4MetCtxBkKRdThVD5D6J9F74k6dIhRu5Qk
e9QpIw0VUQZXD729FGK+MSp4FD/VH4+LndUoYDFDyBVtqZvDY6S8Y5NI5QaMFFSR
XwWvqvW1O4jPdqmf/a+Z6Ps/UOzSS2s4NhWZKt6uaampW3XYJ/Rp9i+N9Q5qpcAx
No43n5MSnIIkm0HGWbPeM2eWGfuCfxuXICqHNn66WtJD/BD+zsidgI7j9IeiALu7
441fYHiKV5CSKCENzDdNKBH/MW+88KMUrsn1IUwGRvTbJivmg34ssubHSEpdpeP2
ZsAzpUKSep0xJDGFHtV0HwtyZNoBNC3tA6D4jkVuA1K/GZhd4WkBp7/TpUjdauTW
6Ii54PjBlqAScNBqRe5FKfPKbRhe7yoMBeDIs8HKLv5SNJSEDZUnnGMcxjZVBpVI
e29HJ65nS6MD3UHLKnJfPltTLUNRDIa5VDT7m3u9XMwM8wJeEL6ahpkbaO97Gu8K
olnUIFqDWT3BOTTGDT/J7T0sXaazn7k5Bf+tgJfctCmKBQcwkQhjVkwxcygyKEq8
bsbz/7V7XvrDK7+8C4SFMYyWWKHJVhPOK+MXeul9/BssrpuUeDxeAc5bS/81tRkF
SBEdTQF/72TBNHAl3uUf992Xfl3DZvj/NXEF50wIGi9sK4adRw6GjC5IvGK9071W
XO8EWwTNWqQGZ12XBtXaJVrKYkb/s/NPTWs3u331pOixQCwPJplwsNUNc2txc7RC
zdlHAw+XRBVLgKqHO+U22oCNugWC8ijhc4MMctA7hxfJ6FGnfA+4ZkeEzXUtxk69
6/FWPPgWgLCA37KyglxnxP4GRyoZIYmumQE4RsyB7dnzKAoun8Z3zlX8vRfWeBbP
0Tmicb8rDn/Sit4sOjXv7jj1HszI77DXF3B14f6pIXuNz5PgrMRv8G77CqN/Sp2C
Locoqgrc/51+wDEUdvxE/titlNkctZTFgjU03qX9ZoxXou6tmyQm2slYJe67nd07
2DDmeYwsGgXkopNxAqPUCsF42Yzpdw+kW55FmXUpbgYQCJqSB64+YBlynzfo3xME
MrbC97avv3GK+78RayFkJidxhiCGsqMC+oOKl1hVMXqE1ifNrErarmMbZECSLqRq
GPbut9G9DtNoKsWzQik5BrIS42nXuSsPIIaF3pQxcVN8G9ciXS3EE6+0ZwTqQzcL
a+vZ6GaUN8tsin8yeAflhSpyVpgg1nzuxjPW9N99RtJifgDZ95XIM3v8CWuQYM4N
DXpSUuO92gIQ8LrquuU4gmbUs7CqtdoH5mg+eU7uNld+Q7uMXU1PoXxGvWpfip8t
qQMvg3/cDxnGDF51ptkEgbt1nuBrxcQPDxKZAGC35eQxTWrurkxCnAN77zjWy+gw
RcQDMptJeKe/Eqg+ryoeXhW8g0DlAbz2V2KqT12zOSdBAQqFxgpJRpTcbU5dHisI
2UyMikeAVt7w5k4SQ3uY3RlRlZPaFK3gz8nrycsJDZRGX9+ZgbUp55yFbP7wX2ho
Ze+SpTc99b/vtz6uTowCHKSV19APRqPz34ksHOB/qITv+jECTro4pboF3ZnJGNKI
fljjxKkzwZ5JyRFzxbhEIhkYwE/dRsRi7PAKnKXj22wyPIhgsPKHeGzo1Z6GbCnv
+acHYR/iQbTfpFkkHiigrTYMezVpJGf9TBop207xZn0mZUG5NhuEeIMSCK0N/hYN
i/U8jsJiKMVJBOAIiCoc+MEW1BQChitceNgGdptMIIPeoX2jQL3ZJ4chOoEAcBBL
/Kbhe4Q7dpvGYQkko8tu+5/XRTPEL+UD3JsHeL+69BBo6ismPrRe7gBUhXbSLGhi
ZQMCUzDWGE5z+4xRjN+wOeLJfi5RqPmM4MvQaeRf3/RnCRkysV8fl4TkRn0L25+A
m5bgtbU4YhnsoMrTO7MhATPhD4XT+O3JOi1y3rtbpa1uX+ADDUrJEX6VE83qf9st
FwARgDZEcWll0H6jvhfx5C3bTggHC3kmLoVvuxa40ONUHFk0CGH7Uy5PYgz8cdYq
OO4yKzNTz+aRdmrHcCcyfLAsBZFraY8WpUxuJReh1Vx6qtwnl98HmwKbcbYLpUdX
1PdUh3kbtP0tavs6cfK5c121sYyNu/AVaRCgK/YCPsa722OSBlwdu/iQfyGZFhna
jhORFW3noEmQiOuUyZ7G5olApmnEI6O2DEoC1KiAof0TO/pNtUwayJvVDFnCKC1D
NIijfu/HWO/rVTJ/E+9Dm3kSyD+9GVz5VDLny9db6s2AfuRwRLTaO+IJsENeKitX
TyZ/bDcbo/GQmgaTXrkkFUwq9Dk2mEYYhzvMi/vt2botYd/4GQ3f6WIeSvwKGUPq
7p3FctgRP3fNu8xfm5NY0GyAx2sekO/vsS4CtTP4j95w4i8b90CyLQCGy6tscUtN
7LvkTJJxCN/CgtbSdoto+nFtzW1PFmDQBSQN5DcW7GWgHnAcK1RuZDPBDxAsV7Gc
5FWETSMIczNcvpNFxUgbkLVBPTG3hFJg15fifR5Mrl7b+MsBIBrdBVmku+Si37ul
Ae7/tJO3RGDtIUXFowy8F2JxSeEN4a57NGX9FIqE81LiBiEj+vEAhUTQPGFdeeKI
NRvCHOvldNMMcXUq5L/UadBcDHE0B+h1NOkYv4nxZ4Qfir2qfphYKKNslONRH8S+
+hl7qpe1ybvdeI7I40w+IhK34Y+YW4yUoMwu1rlpihBlHeFnbGq29lFzPyrc/3Dy
pXa815zKs6p0UfbR+pD3lT15NBHfxIa8MCD8I+whVV4jNnWseuQ+jwZtu7A5ed8F
Rp9cUTo9U/zYvJV2LqtsB/YYC7EOxjoVHNY1+Zv6AtwFL+oBzpNu5z3qJ+fDi99t
RD96qYPv10nEkGtWgmQYhId837FwdLvTFDG49fgyXuMv82zHQQLdJTctIqaqoR0j
yHd+glue3MCd8k684fDrwsCakzxdKt9DXPviyqUoE+9QZAlxPruVG7zNn7YoK4Ex
6FXgPvOBrhRgFEqqWEvDQGBGMXXyYpMWebSvb8vBYvN24P1xSZQ08BNgILlC2sVi
BG/H5PZF8qxmtn0dBxsype4UiSIhQ8hgnOvPDty1ZAbhVB4y9ZwX97zi/MJV19S5
YquCyGwls7roKRMi4hFs79JUZ4g76Iqfp0+UiAFuocTuB29uyTx1izBaqQOOc/aE
zb7ZZzW1FE+T7QYH89ieMYkL97BfXmCt3xFb9vdWCxExfx3Kb1QoAwUEStmPZO4M
eT2no7O0ux+ovvw5Q68IywjWrbpWnxK6e3by9t9H2giV6GAM4fRX58WiMSHMsGMW
GkFhMDi4r1RQLooRAGqzwEnCRN+IXbedzUS/X6eTu6K2KK+4Gus1aY2rwQa4anyD
kOOEfPA+xA9p7jIc12fYsKTm1PFDWl3IBA03mPbwz7jO+x48jEw7/fP9kP66rcvy
eqGx0G9cSgMPJudFvu087A2uFwma7e7kQvWZX+Qq28PNMVcRCOAJ75xmFeQUZ2MO
vVR0libp4WnYqiShqDxeL6/szvnzZUR1rfhRpKGt5JX8bt4gu9ZG2/Av7x7NB4io
bPHLemOfs6wg4raGlxVNz91r93yNVyAgmHWjjrGTS/WHzVuAwR+9O2CUxMZ7smBt
GixEkcruUXY+2Rx2ztwvC0mqGiVrCPwnSjCU2q6QZGlQveqkVQjOBm65JZk+XaNO
BIKg0y7mwUocHSd0f/4sB/3Z3krvKfjA9DR1BeyHIppVDi1vH5kUra32KqoLJKxn
8tczKw/gERj4/ej00nFw40kDCeigPb2JclGV57wiE0N6T9y+yVlTA+uW92cjFb5i
VipdKz9TlF3i7i4h0e7fKV7yFhMq+++CdhjVDbor9vASy5E9azqRbAiqQ4TIxEDC
Ph35UQINocBpxf+g31Qnv13MX/zqXKjx4CG+SFJt9oKks90DlZj5MwhIRXSvJmCw
dtGTNkN12jxRUsHMYiAXZPCjbgatcw+f4FhF5Z7vp7IJeeHYDp/QZ07dIiUB2gfw
eBFJujikW6q2U6IlcX5FrLXAtzoPe/98ud4snLmLcpbQNtTXQAXRL6B1Lz/Jz2Kh
zZ49mHekJeVa3YAj2g9fihVfZjV1d/Df0oAm5KApEw2z5oMfFxjxhJy0aPLanW/f
ttEqFyUC4lBzPAADxC7cyHrZvnsMaJYDmjvdiG15qoEfiUmyAfe7b8GFZxCbgDuC
HKlcH4RPs/9YKAZD/lRg/n2nwY8CW6NRZ7J/Iui48DIii3q0iOta3sJAqx/LOlym
zaHeIP2/mO5xaCwCFbB5HhSkSUZLdLrs4RHdqHfbRUXHlTLkUEtW+AyvrjeA9Ijb
2lO04klyR2aRN2ipzDBljf28q6z01wCUw3ZQGn5dd9bWkwxQrC2e/ETa+IgYlAkn
A+pJK4SOv1wdnASMQWg66hs/wm0nMVqfm+C0MWX4xrzxdQZ50HA5LIcKgjhlRJkv
LmrbSXKC27bkgHQD04ul//l4nGFdplJ3r5q9Nm+xExAIRusukRTeYyOHPOFzbN06
GEYrDcP6BqQrpKdtED20rYIWEX7wfK2BLvYLE2LgcI7mcNjNtnhaNRbQjewgxlwk
WQFXSZTff+hRthGkriXO3/USTSu1MxalGtKy60c3tTC7nVZazXRBI2YhelNM1E2c
aYUgkTI/u9g1RNJ+H9wikH/82NVJSzzo8SxCuqXP6XUJIXcR8FSmO2AaVa42mvut
clxdIq1L+Zt8qXctbnXOVuKFOF3rp6CUoU1CC7s9jVphINSkNIe8nbe/et0IC9l5
4hMmAMPgRwBWbgquPYcPVqH9QB82zRtjcyWp3uSl1kyYYQByHHuQzlO16Gup3+P+
7VipQw6y7HM5kJlVomZNUauyfmIYN6mG1dSsSvV7vOMuWxEGMuzM3AlJX6bhxl2h
3MU1Lf7lUcjLD1UsmTdY/kwcUd/chpSIoqc88+/zfcvrksgufBF0Lbb29Jsf0Ncg
biGdThXgV+XaDcqOErUGQI7xlp9GXFB1omSrJ6hQPiySQSYxqOeYPgIRYpKoStJ2
kBN8cFfUXYXPiz7MN+PDwL9yxLUNR+cVKAat4VHn6+Md+4bCXULjjPwQ9lWUrW8+
qfJ8Sdx+Aq/mI0tjC+njxsEFmbYbc2WobNsud6gyda5acpgeteMgXdPJAdZbAFgh
2TwxarttdA0DPF3AbUm4jxEHA+dBQv0i+zk9iYQmD+jU6uypxvMfCKrMhaa3ASNn
TIlXXGOXmpzQYeWXLUFPM98YtjYcJzR92qK43BE60sHrPTkgq1KwMqAisSW6gi+1
QSblx0oJYYMrk6p7ITVZRsYFJClSeICkoqGAdQT2jz9RDFT8NWNpG5SxdOtz+3xT
KlF9mo6dvzO9trYxCgyHBffy6tE4+8ojLqx6YPT+Hut6Z30flLcjoVlXN/qqZtzf
WL7hjZg4z1O/R1kskO9/H/LJp0GHekB2RrIjKqGvVC7VqGfjncQt3AILm9t0jqKQ
vjGIl3YL5PH6MHUpF+wQpgDwiaV26CEOBMUPv79fCLuU4qLJuAr8Eh0bfFLJKTCg
OG2sO4dbrEiLQC8RpTuoe8qG7KBNDnRtyRDJDCB/Dv7XQKp/NKnvvMSNb50fUjuc
o9ojtk8ooOJiScwVsoFTygVRyZ+r1oTIyqc3VyjyAheKGnsXNJ+1EseW+llpSFO+
86eXQtwpo2BeafHngZ0TNuTltZTVyCfjC50Lz2HAbkslwWongcN/u3V4XGbAkHBI
RSZoBrMqQ5sy1Xhu4gX/lKOBWDyShpBclFXBX0kpqa/goPfjAM4AvI1SBxuw0zoN
vym5zmeJHKq5rIA9rAM1uUacuibYQ7ubFLt5DMl5M8cYCXBoc+Qb+NQS1pOVCOGi
zP3v921h+cEZX0xoCO3+Nys6ia6ngueiwIZOrVIN4DPlRXed/bpyyyNpkrsw1JYo
J8UjarIwZv04+tQsr1NTa0a6QYbMDfF5rFB1Z5Hzv32ktGe/ILb7dPSWSVtXpGFU
5BTAVFTuW7TBp4v8uYSiJk/nd08T3BnsyYs8KO3wYjGe6OX2qLl/4TDJXk/7EI7h
owMU1bSqaE4O1/g4Z6ayq6jfHt2FU1UmhlGLJzOqrGJMhnvDA5GqNkarrgLQuj7z
8Bx+GDg+5f9HtNcZXS9mOlSFD71IBIXM2M66ur3Ao2q4s6/6qx4FxTQHjmzOWx8n
KGiNqhZZ8y+ZXYBe8eU5hWNkV8OZVNSVLPjpihBweYN8dnYwQAHSpKUmoskperGK
NONXEPA4dAY78Fu6BBs+O3GiPD1euRM3V/NGoS+8IrGF0O2j4TLuq9SuCzZV3u4D
MB8PSl13wmRaZsaf5K436uXls17TFIg3nqf8aRba0+yIxwqTGpvDuCJxwzYPnrwE
2bFx1nVONVpNAjMRTTx862iyJLS2n+XihpOcZRs1+3R/PxwtMrkLafXrM073WMDO
h8D2a1jSz3BbjSCxCt4i9b3/L49DWEvI3YQPJ9fXx/TXASULGpZ99cza7o4tOhq3
BxC61n3TzEEMzeSmlPOqGWuASPHDG5KV5kLYTm9mF6BmIoW1NqRItoxPd+F/IlJT
jLLOtOpKsGWt5IWVI+Eqseoc9Tu/QXcCTSTK05PGqIxtRRsiuPLkBdT3ynFbE8f5
Ep1NPc5MXAYVHxV/PALc+dQpPeG9vVk1FhYC6ZBAF7OG12pxQ5AFne06CagD0kJH
OnkMoMoYKL5BrIb3A04uivKQ9+ZhCYcE96L7EaraNa0A0osGI2UXV1vRKE0VN5ZT
+kTR3GeH2Ww6QoK89sDYXhk8cHNLquxB277UwbVSytLmIgJfbwnqombXX1IxWpgX
DahuiZ1hhLsO3Z2Tcl9eFGb8Rj9iifebZE+OoP3eS0B/MtCOHF8HC4QR4JspW+4G
Zxwhwo71nSd2YCcROmXqL3w+p06ZwkhesmCd9dOKepkJTJsgWJ041XgHR8i3WEnc
vuXgtnNZ6AOtKJw3f6ggDsQxqKtYUIYiDZbmm2mdqqB527Oj78UunutyQ0Xx0QpL
QiKbPKw68YlLic6F2GRhZaj+LhToju2XdNpWQ9FcOizkUCCId6NQ8WjDnZVR56B0
28w3lG0JUOtV3GfcCevlnOcoc1xIgjP/cQzVqCy/P9NgUpMqvvBL5TavsiL/EKSB
Q3V7ElR1DMrpbYsajeBKKhbwHtC6OognpL965S0CInZiNu+XUNPblrVSiLm5Llyc
Ngw5MQz9uifE9uB8kbt2xwhSeTzYbtQZJk/Q+1I1tpvzuSFCIBCcHB/nhbAO9hZw
KEU/WJ67l902/We7ZJJ4vGN181EIq2v5aAR91R8XLeVOAHTEPDiblpk9beO7MrDn
7uKCjmPNexYfpvWkxl0uHzzikBCSwMs/QIIQcGNPuwJxws8pBly4hGKhhK8EEc1P
auLU7iwq7wiXRM+dhddP8CpCsTFpYTjCYgd8yV1BHEmqWvxlP58oqRbZJfNltqPp
LcW2wdz7dBAnv3wxlqe/HwXiPGcbqWRCwjMLFkVKs/rM5ICZT1SZv7iDr5/dnd0B
yjQFUIwpH5bziVZdSq56vSeg2PJ3dZFJXm8ESWIl8tiXKqaBSwRRfkNKTBmdst1R
/8/yx9ymQendmiD1VVAPyecnWqwsIaIZe5SO4+AN385bXj4WnQnuJoa8nAqmu/nz
/K1zCxo4SOTQrXg76qSMCIrXe8PCg/SZB0fDgWrYmb4Ct5//z5v4iJMpuk1TLj3j
N2Au4z/Yw89bUeYzf4E1Nh+jVOrfLeoyM7woCQnQIb4K50044VpvPpWNNgK89jkP
4v9c38nDoB0rsKndhxXZCORvQJczls7LTGqvWtXRYGIzYvv42BYKoe1YzKaQo1y8
spKhDkBDljydVTYwPBvbSm48jEO9im38lUJBvGc0878+XIO7FBD8wEVypN0ssoJz
B0YG5t0keoFfVZO5K3EIEmvIV80x6Zobbnhufd6ugiAv/SNwXso3TBUG7/AdbAym
6T9Y1aWNIPeeEb60Os9MWp5OOAkVdX42bnEigiK59kuzYYWy8ELPdqkuGPxAok2p
kQlGphVDTI4szgiVbCJfpb1jlvbYM3lvO/Q4UnAuXQzMf292sO0ek0qsHXfoIBbi
Kuk4n82VLTigMFn9nFplGAZXbUwq2Keg5gvCHqAP4l/uTSQo7i4g9z1Ldd2cJNJm
q2hZqv7WuQDUMRx6+bQGpRX6qGTzTFbtpTRo+EHxxW+ndfV0zPBcxXek9Pd7Su1/
s/5f9eiONR4IG8bwJ3ivnTS9wNpVkOlrbqrtLauGT+bzE9iIQ8n0evR1DlB8JwF4
68rvxIozXoDFsgptqkFiVtbhpKZH4ARHnd+Awo6NcBHx2OPeDBY/d+IFcZkFg9S6
xkwrigNc5BI4KgPyAF+5jX7NPWq/Ckq6YcjQsHxrUJhQpPS1dJRYaQjwXJyM8+yM
30jQJlfCXuOzRlFAimzo5to7TYOQCX5rhYAawdP5P4rkJXxYH9+9VNrNEj5F3Uvi
tsKf+ZQ5hG28LEUAgBtfRS99fBq1fGZBjKNmX08F6p3q5rKFOWRInBhLX0X+1vqf
wEz0XwjavwlPhC5+CUK51ktpAoxIKD48hnIdheObG8iJpPdMoif9Fe1oKJ8R08jA
OQno66N7lm5jebazwGlfiCMs+LflTzfBprSbtqu8chb6ABhhvLXvkE5qm3oa9etu
DCRqd1Mtdx8VmHucdSeAJ7kwbPKNetB0FKheCzS3hzKnAjuLTahGcvO4AMynXJb4
FAW0l+bUE5BA98BuD1XRD26RTYgveuKahiFPAwwPCxQyf/GQ4RmKDBbFz65f1GOz
YfDviPo/DgkHOvcOebtLh/VhaOb9ySGQVqWfTx4gHRJHJD11JSWPlZaYt9J3xlGS
hWeCe87rMy+Y9WlZeisUy/c5xG1qlpmUYdmLEK7oQgP/xKodxuahwOwfdAIvuae7
NdcG9C8BPOszpHwLdl7DvPQwxgRxLcc+lgPm25UrCTz1eF4D+9qUc5gXrV2FOzEA
qAGCSuIq+864p3/f4CFkvY9T7tWn1NEBtuC4jOhN6ovemS7rhAkF/r0eiml9EcXN
D+DwB7w48Oo9yeZJuMPvsbAiqWXUfUWDU2pdhYa+G2PB4SNAFh3AYhtWmXM0FTew
ei5U8LYoMM1uIsh0/X7aWLSnwVibb+N22qFfRzORh/vr5tnyE3mz+n02S0JQw4h9
I0qYvx413V0E5Q0dpVLRzsiATOdPWZxe5R37xsKjVbf58lbhNL8zg6/PlsXD1Opf
BcvlfG0R7cx+o1LVHoPpUb5GrF/iRmeXoKJEzpLKwKvbWBHoCjQvxCoWWjGt3niG
DkSt9FKORaMZlj0W5hBHFEg2SVnl4fWbIug7JgNICfQ7IKCQDMwrTBh5/EndRqKy
3q3W6t9Vate+T199p3qx3u4lKy4t328Q/4kyvsWDN6K0TgJ7VQqGx3h1t2qncyXZ
hRHOOezcJZFrJWxAr6z6VVk+2ySuO44Su/vSajUmxiZ3Ipy/e+vDBidN4Ui3tY2J
uGwpTlQnOQCTaVIMwhSYagJUX/wkaZr8Vt01SX1l7J+FT58miBVWzaFqEme7ZZzo
mZVuswqer+j3JqUUP4F05YZxld06LmYOgfgITEGymSNf9K5jtJXzYX4SWsoH2rVp
3Z0+8GW4C3DlzDCfDtQCCZNnEz4JxpaR2EyvwJDWavQhVuOU3MwAYrBzneYdudBO
eZfgo2llQY81TbwdBemx5ZCflhIiutwoVOXuXNlRsOhFq3DjK5p5x+r+o7jgzLo1
FbLtVNyjCPRTMoW4cc4bG4P3/2Ton/rKI/lyklTv08ubVmVeM5gAE8dFo2y3krz0
6RVun4L4bGT9umO6iQL4iMtJy3COvspSoISMt7WqrLnd2WwG7r75bNPdwr4oTuL9
xGWSpBSscuc6NMjrHjb8ScGX8VixkkQlUBry1d5X92mtqy9t3ARNwMYnZi1vzKJU
rmlo3GOovtlMr7xvvIp+9FBzpd/74Ckhefk9RVGeVRdtIWF1SdLdl0gPHgGJF7F6
IWXyvfHk1ClpbOnKwnos7ayWuEsL064gBWN7lixnDTrNYeW8HFZOBdQ5Aok7EnXr
ndAii+s8JBCDB5JH4rLRBbNGrubkGTnbTOm40e7RnQk82tVMPqT2pPMPUqK/DQWa
DajscWI2+6HJ8vkR0bka/ADTZJvvTsE/MSq1K00KB6V8B67ODVJBHYWTTo4BjH66
1YOY6ybF+gXz6FzmcWPv/O3A8Eqw72KTszA4KS4Oh3WlsYqqnOO0ITs7FE1OV3kx
GjnnUvjpq9u/tRGn/SNJuAqP5uCZzXm6R0oZhrwp5Sd7kfTrdEJ+vlbEgnNOQp8M
ckmJnzTu4D0sFIWr7H12tMSrQAft7kzB/XdzHicOTz24jw52HaOGNuP5/xlYK6qh
dQLKuIDqckrDMj8TLWF5WBnE5iAh2RMNfRv09zsWYxBmVHIkF0RwMZyiGOCQ4YUl
C6OijR+IUK46bDZ/JyrQeiKgpY1LEHvvaVAV/G33CCoy89UU72rZu8uTtXFYip6w
MNn2gPQpEuzuE9q55cA7DGRIau2AzwHenZ/ugaplntar2DbXXaqqZ1aBk02ILZLZ
81hokvoYvcQ7BLiBTonoEBv19UwoQtBFqULkjGK0YJ3RMIaHOhVK77S0qWX6N+8z
yX0qDf92ishtOvre2Q8/mLNaBmJoLL1JtLZ1fCYWnfrKEFhVFZln//Xnrl+j+795
Pjdc1TXIq46DXpDcKAok9wSnFie6UEr5VsLU4M0WPIwDR+hSRZzyW+MkVjpwcxeS
ocapIRMgObuM/mx048jhZYZ/e514TVI7WQuUsomAoYpxn736tc2+NVKCgmFvofJ7
APyfc0D0Uta2i0bbhqpCCdNjsGDL3xwSz7UzLhJSRntLwKzDVhgXiOKHSqD1nsvW
FAKOdTQ8LypebNU7wJ1x2wPSL+MDj91V5WkdbrYNcIzLyjB0Q/Puhr95vLRZwTTd
KswpLabnlUeHCWrBPlj38nn5j6c8LD0ag9yHHJUTwDNQrXH+I8pc7DoWCM+EY7RK
Fv+Og/GWw2x+VoiOQoyItpPLRdKKB09uEYD3xSq4UcqQxoJsOT6eV6ajYMFdhi3D
H2cVupQ8MUXDChFVxqat00AEe2kQXSsjZt3ltQcEh2PstOaloNUpc91rgvuZ/KAa
ETm3nBjb2GONZ0CWhzane23cq/yD3B4xFwqbTdPJzorZugl6c9FoCt+H1o71dx+Q
bo1se+YugONhQrhPKY/2blDI0wHX2tTzcxfLg7QV8OUGd4j1wNs6b6A/akhqPpLb
GljQzCFbP3Q7RqOAYQohxDikuGqwhPBJYlx8WGhmz9d57LFc1A3nv78F7itDxRuO
XnA5bFPtQa7nBVbaAP1WEczL89FLBc/bgB08o7KwgEVZtuQGf4q7jlpUW0RWvbjn
uKgP8uaVl1kjycIYEf0O4kuOEKGvR1Wa6bxmPtBQ4w/BGRPXFeVnb+qetgelEVXi
6MRU7A6M7Iwh81RX3yh9Uip2BHnp70+VLWXcQeknlMnGhWU6AA2vGuMpJHuImAr/
nBHoFvPhAT3D3q0+Nm0RQBRnO8oxcflgGM/2aqbgAkD/PaZLz25EOxHr+IKD/PNH
F4KvpkgZup4dE4Kv3zWMn+umdChxKJDUX8Z+KUiEN2QiPkuzhz7bKtq5ESm1ynqe
2skmqDMXgjCpuauSTmKCT4Y234wV00oBvzKxw6voP+DVS+YcWeyS/gJ5niYY0ACK
aC0VXArNWuUp6GZb7m2NaN7TsgX49QhSj0kzX2/SkQYy9o7ckQBptrM4bsCAgN9X
eL/3xpchAo1dSyupZzoKwszgsSynEw5ifcNzjDDuIrGw3vj31fkjCDV7fpVcAX9+
TvWN2/3qILl3WX909k5RBiacwxjfZJajcT/i3FVAzp+wpXzhTCi+67T3x0xz3ri0
JHWAroj08NTcKK+8DsENB+MMAUOMbfbQWT/08Apxp7aVk56+oLfbyeuawNASJauc
Y0p24sVRBBDs7ZfSDpT3EJFMhySUgiJsTMT3b5u84TZDCOS5OEJIR/uKIRxkP1FR
JSFahZ4LEh+V77I0NDE+JCcpHCG/31AIJPIVwwsk+txcTpRYbiwPFF3bR5QVazCo
2hm1FlLzJLhDZE53aB0Rw4pkHMAkY5zr3q0N7Qp/oCZ6YWIIT6cQHCyv8hULXoFY
joGetHj5i5SxPxGQRdv1hJbmiUwNVHJhjpukfJ/Q2aZlBb1lkzLxOXmtoq6pRAWE
wkrUb/rkpcolsKMjQPZdWtrtEFjlOyv/UeplwB4ebZM5yArPwOc8/spNDcYa314s
shd5eUWvMVfo34MLCAUiwlJZPCxDrPlyBHe65X1Egoo7JDip01ErPewyCbodxHsf
xRhQAIwk3HVDD8BnvCl6ZbY+U1AW62HbF5GCYgDu4UU6fljuOp6F9IozJxPyxEaP
2J+C65rhIjRqOuCO25JJeTcU/utG12EhqY7+SiP5ZTklUJRy7sF41X1lz39vgIlL
3Xp5AupHm2t7cyS+2pZyGPfovcGO1/QC1nZ49ZyJUUoGw8c5YfhukG65tyOEQTbs
8eGgRs9+nQ8U6VA0MXsy4l4ZZu/h5bY4TALH46L0dEMHalaQJQ8+cNJg282wneXX
5L0hcomR6uFcbZ+J6+Wp6ITI1L/G33psOuaPaq6Hhly3jZoKn71PJZdy0xrMoOPI
YcHjQBVnavI7XmfGBIA62fi4hxs3Xz8Jf1Ujf/eN3/Mn0BW4+s02QGoLQIcfr+jb
mOpiJds3TLRUY1b1IE7gUAsSlg/7bVecvy8GHTUGBlOLMi4eQl1rQilsjCoInMfW
gNvNv7q3tfh5r1NI7jLgijyqbLpH8De2mm9F1XE8h2XRD46VA3Nry4+ViUS6xRms
JBkayX92zSOKk7MebPZRo9k5q5mIXOZwxr5BLmSbndIl1/MeRkPvWMD3eS1uNd09
Bxm3M8mbev56jhfW9QlSi3mo1XrNUjsaPcARgNAQXi0py0oDjd15dAqGK4nweAyF
e1dGgZ6tGC9Bl8nAEuH+6twTVviCkjxt9uK0Nop7h1ANYZxItyaJRicgJ/JH8Xak
XN7bwWqCmmno3sXWQ585WYMMr/VWke6A2tOnqL8vjCD1XRhGPiSAKHmXlROBnm44
Z8pGym7uRYq9PDd+LrLOW/2IdDW2hnfWGSf5XdHjRcbgQKOLxsme65Z98fnvDJFO
XVp8SLExqJNulhl71GJQ9FDG1BuA3cXH45t+NmshsjmZFEi3Sk3x9p918jn0g4Ms
YIOoAQvW8xvpzvNy37+ffIIicPsPH5NBu+nHsHVyTeXx70kwKDkqGCh3LNGAyI2D
XTFF+reE2MDPqjw3Pqm11qAWAatIXxx5q/rjjAGmKWOWHL5gy6Izr7HNghrgjWca
aMF9+jF/TCKLwk2SYEAzqxh+tfIUrTBA/ZSspK0yEbCt8K2EROzLM+SLP2R0asvF
HCd2gvT5tzGNbVPC62Pvkl40gkkhAJzYgDUsNAgnRjpviO3Y+RXlwkdxB/7T5tUs
EUMUGwbt1NU30SjHFYr0nrlT+DN7/cHNZPccTs1/xLQ2U1JDfNnjGZG+q+0SlMgj
k1M9MuE08SuY7uOZ2JnzrCtNzhyza7FuGQMYJNDVpqPXdcFAqB7SdCKebXCxrVhM
MQPUmhLjgD7rOYjPpfrnKS9KtcRffMjUhSQzt28lDzKPrtKM0JJyEK7AKiaa7NHM
YNWEDDxDlJYUHypSMiDdEmyxY0JE9g5Uj+F+3RYcAIlYGYSXFsNQQUKlDeCQfxEC
DBH5+YQeEmHoyJtfJHOuQZlcrTca4ZdvnFCTEJSNsj5HLzlmgEKTa92D8fu1EWlm
EGKsVlMNHRmj7uEnnJ3SGCdRgY1yftfwW0w2FegziceRyT2Mjk9x6QsHNAFogSYa
bZHacm+Drd0UTn/8/mFJdVKYtz3bbpsSDgZidpJw1q8e+uMDDILmkOO02c+30IBn
I4HeEX/caZ1ujhBgQ0GDRX4jm3O9VMKp9boChR6oCA4rGoHry2gFMlUEOcbCKxxd
vp03RN4K2gudQ9oLEKmmwxroHx4Rd16IA3d4A/aUM+Fz6+zL7mENJ6lPP702G0PU
72GjHbcKwHJtTPkvExmXw+lK3b5N4A1DZRlap40w6bZgXUbTe7JiL+4xbI2DvIFj
CQrnQWXzcRq1mGaZ2a+UTA2nheCEQtPABGtDfAsYqBY65PLXJncZdr8QPJgpaJl4
6isklBf3S0ZarUyo8GlhQ7WvEdib9Gp59LGDJio3IV9vyfBc3rWPpKOrsudtZb6d
H79w8OMujFaGRpiC38Odl5HtkTPLIvrTRaFVG6h8tdRqPE/G24GjaTkqVS0XtfaX
N9FKC6CH8qIJ28wBscGBA1fFnSGszUbL1Mh8K0Az93dM32T6AqioK+psHHXi/Jr4
NgSpNJ52G8gW6r9xiLScPUfYGI24yJDYZFoK98ey2xxgJR8oysJAJhEWkICFtUCt
md/3u5aFMTmL03+mqHQMtzGIgPKUkLWJz540cPDn3usVcIs8IScbS/pEeLLogx0r
NgDEGBQt0XNe6pfgxMoT3cWXvqtQByl3iU/LOaqYi4/6vo61/GPkmHU95oo1x+ht
6VKz26jEHAOYo0XTzcYrHtfPPNieNy0TxH0LMlvRlEY1ka2RB4sZH520Tl14Boqc
RzwYmI6xvpFM9qgg2VIhBQODfuvi1aRINKXAATk5o/KjYC1JsSpX8UixDTXrH1Fh
fCBM3MeBX0fxfviCPto02yEwSYI0iu1uBskUOgCHgvQQgtrDXwvqv6qxi4W+2sl5
uAu1lFNvGDt1IxJMTsCMQhKjZ4SbA8AUoDbtpyneMuzxXxsoT8z9XoglzqwfqB6F
jzVqYVp4JK9hTsopgR730Oyg7ZeYMjccxtHWqO4gDhvHicH0+/RV9Z9HfQugdjy1
HeDVw2mom7PHi/ND16VBYsYKYgfDxk2gJR0L75BPuc7f+8DmIIh54J/VyH3zSAxk
EeVtClm3yXU+2vcB1m1T/EbkPQbCYL41Si/+w+YAfyK6KnaL0cCKXlTQGASkHb0F
3e9Ji0sS8vdlXyqf19YbgWOA13YO7pssdv2JB5lcYtvf8yIrxHNlpRVE9YR2CWlv
jw43kNg9sgueOEHE0ERlHy+4MWD0yz0Oj1c7A8WX/wJYgkjLgPau8aq76YP5g72c
LMP/8BsnrDH7JCYxVRPNKJoXGrTrqzcPKuZB0sdHLhDp5eaeJSGw+t5Ciy8g1GHz
ELz0/RUTqeR9A8NAXSt32HPz68FQHaog0nGAy4SYl61gGA0OSid6nDm2TFdEkWDr
2G2d35N3oF6eRiGNCVyM8DgM710u1KvWV+Gk/JYFppY7+VmZ2v6NTdvFDuwDvcFB
RjGquEGgKPPXB0lCgRnrsF+zPq17AwAS/RiulfkiVfK/0AxfnzUz2W9vUHdDeo/a
iZpFrjXGAWFxqdQWZWgYOB6tRbohyO0lhJ3257K0gMBkNXeMoMU7/tSIL6ZVS7So
Vx4yiNpi65KOQqi68WMV1rz3tIrkFrlABfO6Cr0wV+kvgLcweSVMnphdal04B0Ng
RGklg6f5flwmfUFWXMeCn+bOTFk1TJLQFD/SNdugGdz2sqp0Qgb9w0LLJKagKw8j
BNciMb6GaxNU4u9b2P9YXPDfanQsIwnpV5og/9T+v5SfDRBeOjVC49k4PY85rQ5L
gw0f6eedk/4ckxFxgccGEY5LOVfkJlSe95hCMAih0O44MnMwwuDDljLp/e8kwuFY
dhCyJOB2N0uhg2bctbtEl4qjYetDPPrunGbAkHG+C5ul38evlOK5XzglVWdven1O
FXxaGKBpx9u2KoTlvItlGpJPwU29fTaJbdJTDNTy25gWUgG7w+Gwt9lLoYwC5D4w
oBdqQmwhgDY0FGOJFyZCBAXvaYDz0fAl7IE5BgP3lnPa+gwrYOkdHdkq63KOLXJ1
j5IDmRJXnahAznGqR6EHmdqxJF41cjuSiQid484aD2jN5c5BpT3smhAH6ZHMveFq
SoG2qq15pflPSj9H8Rv0AnSBido89i5xDuZAeCYAWnKxLZaB0BtTN8sKDmY/a/Yq
DffvVYawvuWySjwW0NLLsEORO7/vJ/V34T2UQgp9mRsW5O0GCWS47sgY3enSssbm
18wog7MBq9I/szuJc2+nv1f4jhUjveJ1/Ri9tnKiWGc69WlfnTnsvePRJTRGvSPE
X/RNKbWNEU1sitR8UeysSk7NPQm4MV0ggcMmj48KhwBqxUdL1VTpAUSIkQaWrVc/
zcEYR5M2zwz7DJyoavY8IjrljdbnuTcA8uGDnWnOVA2mWXIgnqMPGIH7J96m+toL
sgRywrY4wtGyy+Z63cPIz8wcTK89BxBNxL0fXnHiQF+dbmr+jYuW6BgdNcxVptyH
h/J6bU47o8H/Fe5hMaUEYrj4eZgiivJ3suEtthrdwRhZgMW1o7LPQgYZStHVtArJ
ErXAp0ydaVo8Eb5G51fC+sHVOv1odlTxMHAdMuT1S8JEtMu6vLog5Ks5vQtM+vhU
3Q2z0SYR1zJeCoM82DoSQ0K1vYxJ6hbtnKGh7uvbfZoLVcpADvpKMPYJx+jO7CkN
F3TgXRqBMHhPDHsRDdcHffq6BXa2QKgQlTpkJ1NmjvpmmTFDo9ObnTyXQy3HIqm2
cf8Egc51n3UfrOjyOsLI4TgvDyKywR0Mvr6BwnmwdNI3itYhxtP5D3vSoUNVHqRw
XHCxX5+plvX/xWqfPTBi/bUXB+D42jhkKWNW9wcvfgiM9w0fREundL5CXi7zSC2w
A0fy/ABVM6EitE2vaEoXcx/3HQerPehRCE8sjIpBsjHclI/Wi0qw9mkkiO243nkY
1C56ZnNWD17uZRqMosJYcVzWflM0FwdIQk2fm9qysrRf48XchDe96qSIAtv+FlvU
z3+7QdIB5W5dTga/rQGux26/sxTKTC4jWJPJOYXDhJtEcFaE/m343wB47359gHhJ
dX6R9DgGEC6v3DMBYRqms5Kc/pE/sQBK/WPwx3xIck2X79edASiQaG0zMR0ss06V
aEovu3MCUqq1sHsrSg8REgfWvL956YuE0uQN1Fy9XXvcq/jmlRbnSuTg+8PqB4QE
CvO9+bFUvyx6kjXarxHJLm9poI0RwUV+IAdsM54SNcPvoy2SL87bxMLouiq8idYt
qaVtzUE8v/0EfD8LUJtwZe5mGd5+1Q/2xBQjFpwfu8DZNfEoykreX3PRvcQfYBpx
vRhMMui+cOKKozxyWr5NyIvwB+9Q35WuIcOTgLXHCKECnj+Rb9rBGrNBIzKxfcFi
2rYVmqi08cEHjr0HLBhLjzOHqdgTwGlZfRL+LpD8A8qGL9SgB1sthlmn0o0LnuxO
8Wni1ulWMbQXdRy4wwH7DmKxStNOkWYgoI2dtxXc6oBZZW/ZLHRt5BS/nTvGCHor
NgvfmkzTQ4f7fGbFeIJf/RRTOPxU4IMa93x5Q0L9zH5ZZ31NndPitVlR9F12iM45
i7sF8DXBJY9O8dofoUxoFZKxP3p81uv4mq0Hk7B6w2UNRqOO/MYY9ucGx4ZhsogF
utH37GHxs8vtv495yrLQJiuKyFCgxiUOcD+JTEHfPKVXC1CHaMIDCfnEYoScMNjf
O0aH06tENGj5+jkkh5UpmMTszKnAvpL4OzKkSr6T8ixfM1L7vAlRZwTNqTmhpqMe
nHPMlfTtusRWzRg77WFFQCgCrD44KhK0D/IVQG1yBW0iB9u7NW2m6ulk8sxBbSWT
/2ZrXcNw2jX1EnnrBLBT232e4v5HJdm4wEfttbyMjiZ9leqbsEPpDLzo2X7Ns0NP
fY90XndJU35rmgLT2sfyDZaQ/Bmp+PH1mXwNHcjc0bbAN0JYa2vAI8PX7NSU69E+
RycGDhROzkbs4Rw9vFUsesw/jp+6nK2033F70sIMDvlLxxy+mjQvub7tG/eJPP3b
xW5iUqueeneNtXWLYYEEP171KUGR41Ci5R601TV4Awnc1vJd1f0koeFVD7DYwGc8
/I91lQQCNBy2mlzX0SlIWAS2Zvcy0T3HO2vbRwx+ewAZAroALA3YsL/9yR/sWdkf
sBFZoDNQIWeeVQGdn5tKIPB5ECU/6WyLpFkfi2x/oSiAkoGc8JvjUfLREJxPFjTo
9XL3OxSGfWVA4JBf1ZzlAqVrBiEWoOUGIdmVBElTYxQpwiAQUis1SmVpAw06Bx30
hJAN+nFo1ra3Ai5NseLVA5mCrFSH9E22Kwsa163X6b5pBw1rzTq12/pemktsSTD2
kwSsveePBhxQc8CObYjSSvC949pdISHaOGiJUX+b9WNf1Y07LsKbqZtZhwz17iFv
8Df55WKn9LZyDIs3fKl1EKSKfUJqxKQY/HF8Xp9/tlNrBvUvbw73Oy36JW8bV9iA
aG7JHk1KESeyTljGKofUBwIYMSWW3d9vSGJepme4Yx7ehHAQf7UA2Zh5ur/wY+DA
YPcSM1C+l4sJksuRV7jxDGDM/Ndzm1XIZA6HnDESKkIYdMXxRsX2y78DSSFYrQl2
y2rv1KNytAThg7iEXZdRBxtWk+kj3Hhqu045U/zvteGGlMZonWjXQ10ASz00kvw0
MAFqHB6DWsj7i47FMVLBlQLV8lhAToK660E99Ma/kRbQncAkmQPVErKL9gpjTe0P
/4BwAF2PH0wbfkYnuEz/mx30B7dyo4DyGfDtgno0Ui7aH44RJZQumGKgSDllHp6L
IRCXPxqYsONBQSg4zC6V7MIlLkV7m9SbrmR9GCcShnkl5e1WyOvXKF3K5ZeAE1lu
1q8u4ijn9AZq5ml7CtToU6u2zahFeAbuuQ0hLEZBsTRWflzThtfNQmjN8RpNAA8Y
AK3TcDKcDIyq1+oDeNMX5fH5+re/8Ghp0oyc9r1XOVshQOqKcYpUb7/hJ+IRXv4N
tXjA9w3uv49VTL2GKunfRbiKYah/68qkeYCNcfqAYm18x0LHykwMek00b8IhqeNU
+xWF5ez+dMaTlI4kuMYhE2oEh7CHa1L+X4T6s0VZJLLCDIHNfsiqD/XU/uZ8iv5E
/eoUjjKMW8LQkq7wV1ckCcICT+To2RXk4kNuYNB9xo2anYlY3+3WgKPL4ufRNanO
EvtSiAP0WQsso5B4xqOZDZjP/rh8nYbqOuTRxWA/kywQMuNpjaSMwj4dST9rMKVz
mGMXc6MWI9sZEnvGAQ7bMW1kbMoeOfiGenshMguQbDgvDOiRvvjvzOopETC9kCNR
UBrJ2Jqkd1ByhUeVjcVl+YdmLH/pAvS1pTzrkgWWw9zKHFyw07kf+vfwnHMnC+EO
GpjfoPywmVLlM3ReWKFuVdXkKa0s4RNhk0F0bdwivkqDdvFh6KnB+D/bWZeui/Qu
DpwlTQvJB9jidvsv+T4zfCy9JuLF1R3ArrmIRFsQ3PxNoIOliQWp14rOH8wAQ9qz
zSW0o7Cr+fkvngRoKM4WQtcn5Mykj+hmwTiOrpfTDcJ1kJK6zieSQKS7tq45g+2n
CQU7rFZZiMfoQzvpuRyKmJgkFETC8GTJF728CODrm3+YbzLARUdHCRtcjCtx3T3e
ZCU8IvciJGnE5+iWTn5Srl85cdfeIcSBasr136foDf7dQEQqH2Bz2obuMY6umMVF
+gbbg610DDGJVwY1lOc0EsAXjibM9GveTc2GqawVDpa0/AkW5HgG0OL7vU3Neh5U
+88RliULlwS/G4f+ZCdY7i2IUafax9+4CPTeoqeA2p6audApcGJ0eCtFFTVZobxE
V7eSRj6/7G1dH8YrSBuMQOHnPXx7+e3C8JlzzUv7v3RalRxXylL49upMhrx7vxGU
l12Jma/0ZvvOqTojsdEy2NbRtGHIJ9NlGZvFIyx+kop6aaqX1HLDLSb/XKR01/6N
Q1ARNQ5j0vc6d0rfDbngx0vEMvdPJkrpLIntL3ZEnirzgCimpqyG8GntrgBMHo1A
erldwZXXvQC9KSzkxe5ew/v7yzTCEoRmRFcKfFilRkWKDGCOoqI++mxNRQ8FZGFY
2nu0QRqDuu2Nf/sYqeWWga/Hs8ZtidCg5kodhb2sGXHEsbdk9lMu7lIDTtma3KJF
nU4gPgQxdHGVLvBJM9NApeVm0ssVumPfq0enHEVwkhKcUUBziHj4ze/lSJwZmoNF
/YEKYbHRymnJqsY33kXK2AmRPIyEajndeIg1415c5Xq5fIp9NoybMmfkudCABKLL
G5L/WgrmbegyfUL9mcXCWXJ8N8cbPDHpnN/q3XjIN2DyNQEx6WID7DSK6HYMHQiJ
0q0ikWf9FrzgGIDTSgoX+OhlGjAhKtFluGRN5IK0iH9quhOKFnQTblwrrQWtgh6N
8RUaQKdWfExNkwX+X4fhTox90a9iyPSTeRA9ZO5GZJ0flG/aFGDnkGraYQm3y07f
Vq73HJWrbaOisjpcGpEYbdFtrsqxJTrgSd+zMzM0YqbD3kpzBD+Hrha2HGSj90t2
3SlM46/hkESENcWcPCuyuHbnA6UoSDTkV+jBT2A7RzbA+RxfHzYgssBQ4IcQNdqC
EKZlCmfr4ZmAlGHr+S8d+S96OVq0gahhbi3XLiPZ3ErL7Hbe7P9Je21XZEyIPyxH
4Jvh8MIRkpauzGnFLkqu73HQZbS+eXJTNSbVs4PXzyGFKyWP7j9eVCDHv+3kwTew
cZYoj/zfN2cNeQUEoxMTJhD7Oxa9G67rk+62pJfzFlP8OcpDPb6k3Yg3lDms/M9x
GY+2RjwQtbH0XRi+x+FUaSnycQDyj9tS0Pj6HxNGZabKABU/iSOQvVHsjqt7sNIZ
AhhXPNXP0/zSuvICxLUbMs5r+mba8UJYtUZ5M9MmU0/7Pu3IeQnokXxxxoAPYCPL
AKFfNkkBlF0I37OvfBhPAetxmxXEo6+Re1CY3pwPEcmxVEuQ+IhXPUnhFiZ/Bw8Q
t/JBViEVyCt7L76HQbmy9Xr1nIbIN1D90ySrrv/zqTK8P2QakSFZq4ga7UhLYCI0
gsIC/5gCyoYjuFEDUakSnTz6ALtUzSvqx0/oBwj7Ba3ebATr93iZmPaEagEYcqY/
OaPE3Y1OYqHf7NFXUDz/KKcsBhXDo+f5Ow1p39lkkzXpff8TFsget96iI32gsehA
v4taVr/xNAQS6e1iYn9M7c6qI50sslkmi04ajgGHXAjNfoGb1mi0+Wjrj5Msy8Ry
lGp/SocPvg9rJBHzPMOq/c/ZiUMj/o4l007Twk/u2eSSA9QS1+qAVTnPVtLKPmjk
6xlC7EQnbmKI4jqpR5MwjbkKe+vhzGM9CV1Njm+DygGsjV+k+Ps4qFoowUhDEIsw
KQrZuH5+T24QtQQJEWmgKhmxsa8b0Fs+P3ZEuCFV9h9XN6olZrndcNKm7AbmIC9U
MOYn5bLnvODnFmfpSq1Ckr7TzzYDiU9q46UEaQkgN5lgrsaXoMtKspdNXLVfxNgy
nclpIARFV9WXUShndUs8ZN6L1VsH8jiVyFCTuHU70llVTebDdKmDT+EiX+GT5Td4
LMs9FFKCypWtmOZoPlgUGkoy+cT8U54U6DvuqFQlrtYhnK3JXJMtz22aNo3xEwjX
mhHIQPRdd3njqqyFcRbMcODAlvAwoDsg0aKzuk30BaTKk1eYRW90T/Rms1FpwuSl
KA9RRiMLqmQvNjLFXK78D7zVZCF0+X2Eh7J4RvgVA4UK9Brrsp8sSnS3eDEHbkRE
8toSvifmwoX2tb2JiV3s3oxK+a2bOhUMTXLAEjuG9e+9dMczVOxIW6dnVuf7f/QB
1yTKu2rNiLueNubR7pg16zPAthKqm2BLvxU7woVu4ZG9L5fRYCRVwOEmve7VZdbh
VbC12vEy1phTtCzdmLbLJ0VK4AOFQZT0YVpPaAIXjtiIpMulljXpS51b4B8Brytb
vpNrXbMHLY5+9SAyntdGxaoMs0L5WU7Het8TbWCuarUSKhRPbf+TnyuZt0qG0mkG
/gVQBQHE8Prz7YGjBB7muWxJLOw3E+eMIWrAzk/iU75Ssan7MvwnsKEl5LtqpsWd
wrW3YXGOV01gx6TBKW667VoQ+mZ3N+k0KFHKxvYukTsID1tNbthyqxSOUG2aIPtf
VMunNixZbwihVqJgshLa/suXTQcHH+7jb+nhU7B1k7OMiqDH/C3xKIcZ5Yd5aHaP
n4AGaWvK9zKHBE9Qr4/rH2OnUmHwHQWAbKPTKPIM26usLWdOtxZi4KJzyRVmfP1m
jtYGwEZMCr2j1FRGRY4Gb0FSwmvtUaTahIYmsLFjYdLFT90//DXwFWv8bQ0w1uGS
N5gLbefJHvhbtKU+1POaKsxkwzAoQwznOnJ98d9diU58pJ7ockLmDOqLTA9X3ypi
hNwjswYTFPr0lgvo1XOYy7MCWg/8K0hq3TZieIZZ1ELh7j/I6JMgdmUNdi9Z22sK
aqMs2a22PMyqN80PRbqiKZpKbaN50V8QSGZBbflyvwI2mR/WHuTj82iOFcOrjxGs
PvZEwkt+Ic5b2ioCIhtP5fqK/yJJQIj+gmy5TW/5u4RY31lfZ/6eCONnD9BZm4VU
XOwPPAli9la7v0od3Zh25MdbBz/U6rSdrrsPWKIf8awF/5wg62CE3zIyK/exY9Zo
+oUmjCRI0d9XUtwdeTEdwIlwspvi86S1M1DPHhBx8FRpi4ctkLJQIetMqj3suJiP
eAozVf/+qMI6kbElstK4sqiJOYHRdQsnqPpuQTKAbyyGm6Qn1klF8jSc7Tl0zbP/
Av7QqmPa+MLQlAanS+MLXTOJJxVqcqmAMVC1X163ITakoQUMgMUqIAoR5YD5+sWg
1NsNtmZRLqUdHtjzB1SlxoXGxFPAxJ6RjcnBFKRZVrTtaHXxMqLeLYDF3GM+VDNz
q6Y9bx1NqC+lPD/WW7CSGD/FUflB5u2lUxX1ZPwcH6ahzJZvxuKVTKSyElntLdtT
SANrbx2PllED2XOdHS9CB4wk6yrBhMt81zffDxfdYkmw365LA+gis9VTvm1Mjp5Z
NJriBUfke7m8FHHewNT0ycs7lpBdYA1LqZxs88UpPizdSEfGOEpNW6mlccJNwRDu
x/ollkIasnyx+2cLHl3CEvWkIeYW80rFVmI0BY0NdHIv2zAEWUPq4YZBmKxdP1l6
hhhfTzbeCHEHRHTooZzfxJ5M9ZewBAQ5WsU5SXBSoS5RUcxlUe7rtS8JmPKSk81L
7LN6P0Ksfu1jkMzww6a/t4nLuYfYTlYqcGFDsC7AHrCLDbsNl84GkBw1coHRDZh5
b3baVwspFAc9ohQD0fN15y7kn93dsOT38uTSFnfJkYQKpjIWk9lMpPRUoWu4JyL5
J2OudZh4tRMjC/cGYFb0pRVK6JYNUWrfG3rS01JB3EWRWI2a6GOmygJelneVqES2
688bIgr280czTlF/xQkG5GzYq5XCqoJ98LHi7sPBP/2dlH0AzjMZ1SbzxXQM0ikh
vupmQNOURlnDU/xrKSiCQe662BfYFcJ+Pq2H7HbVRfxIhm+8mz+CVTjakagRWaC1
58a79Art7O7S+UXb0W9+GnUjnQJflzHlQpyVMxbvjxTBLLD+IhczDYqByXIqVxXi
m5lwgLP0wm6d7Cp50fvZ6ck2U2cVSM1kXSt+pRF6U/xTFAPePE/8QwUjBknWEvIs
8w56XaIBcvmIEgu7CGYOBbNDAJEaiM6cjTYo5P9H6MKRqticbcKZ6YlXV4cJ2Zv7
15tF4PN55D10jdlEybN6f6nNzIy3k/FPzUgHvP4lUs8H182HsYx+/pl8Y55KDwM5
owy6QY8EEWo9h9EXZphMVurFyKYFlvbr2LhGMWai4/hj3JC49A1NkGib1feOxNSa
44jVKepqRLJqKnfod7GMVjB7J3jCz9EF3+Bb4oaAvPmbroQakYuu5YKpdeClJs4f
U5qhiucr4fViD3JHen6p83aC+cnNqCyeKklt/5JOfLEV52FGkQm8MNU/EXADIfrv
Z43a+uJJ6fzuwlxDZDxdMZL9p0GyVd8hXGiRGKdHAikZIMC93XEMsWWUKFhOJ0G4
zQlESRuQPZR4o4ERUgGHcL24I5a9hrWhT1O6eMdyL47SiqBBspEFXpmQe3mJjreF
XIr+iA1AWdfy2PMKtI/2BML5UqFVRgOf/ET6cIo1BQre5dODAnwUgAgfF1zky7Hn
lMgE4Xr/Gb35PyP8Fo8gTRbmIqtrut4vyuu7F7pfvzHHItBEATv/ezFigVuTPPHk
2u+gK9FQKJSqDmO1g8GFry8xYIEVdWQkUh52D+MCku8sepJeEXJV+BpqUvy5DiCF
fPw8+oE6vA54K/wkzzF3YtLY1ZaxS076M5F5dc0HYW2wGXCAzOYoJOT4NsjtFYFq
jtiHqs/AA7r/GTF7asyxrauDT0RFNKala3EZozyL6YK6+rFbEGGhWtBHEjh49xpm
0KydkB3BoxguVMwZmh/4kmZHezbDnGxYaeEylprgFWlnUh/rrmws+Y+VSsCY+n8S
b5GyurFHzXjzIjFlSSz/uafO27fSy7hg3R/7xzCYZfcoCexsUr0WbOSbVmWiKXnh
K9Ahju9koexSCqygYIP3WpJcSapboKFfp0NBTwtTtCzVqpVKE092yJKeQSXizNbV
OBigR66KYmiQCE2fa475GUAuKS6VP09Hf3FaWr7KSX7wyf8UJTrFRDR0DWb+gZl3
Q78DiSF3OLhEQL73lpBqKThbE/DYXjYHCORfdeNPsjHPduGf475b5gn+L8J/oDBg
mppL099kFrUhkkezLYZmWGKho0OFSfXKREd6tVziyzxLxxrzJ3I2Q/Gz2w1OGpA+
0zHByaDxWnlJY+2kG+gTtV2AnXR/MqR8T+OoDk0gaj93glyYdNbskkWtVbx63xKr
GrWggcx/Cacu5vaF8EqN3BVxcwqUooH6ymN3mo+lMtLuBw0HNSfUBPWiJj++tuTg
bqbAJlx/iNYLR7y2PjyWLJPEc0P1NK8Xg0+HcLLe6avb/TXpkQKGs9CNBjCB+UA0
lJDBRIBUHRt0c+XtvCanf3SVZmmw1oPBE1T/AeX0wlb3ElNPUajHfkXxWREMAKqH
+xhf2DDWwMXiv04QknHn8HlZdLFjO/zZEceHdGNCM9fRXox55Ls84kVB/gH/kMke
MAbgIPzrmr2fZdu6K2omIR6dJs0kQa8gmGqyZgMyQFB4P6gld0mTCXWai/FC2WCl
1epYiik4dmTpJkI+t5UKx1kfgDzpBkk7e7Y+XJ3kOFqalFTD/DNMa463iOKe+2io
YdcjVelHkY2cF4lF/2vUdn1w0E49KZpJ0OP/9n5Kfn8yVpjeiwssyVNtPuK/IQUx
ri3zHfGXKRMCkJ+zvgMyYbTjPue5EVc2+nebAkQN3bVUBmHKSSFYH1n6LYRNN+xl
rOwVq+Zv/fKWfyDchNi0RyiCQij8dnbYrX6e01bB61uSraT1d0i/kK0em3xMihac
9WOX88+16MMAUzBkwOvJMAGOK7J6vPxvjWDoChZJ8AGdjaNWdBLQfpLYN8YG4fU3
Gqux62dCZRpjhTAcNy1C+Vq5/kYAMRjFkU1tiR5rwGvJ7UkTQ8LuRwSFIY/PJjPs
Zn9lvzZb8JGLyidRAGZ/3r7LWBC4anY2FTq+R0HgoOmHMffXXqS9vssJdwvuEQX5
Hq8Q2RfGpEO6iBUnKRMZoVqqOM/DahJC7Yc673wlxtITJ42ynEo5irzTM/f1+49X
BIZogXPvfuwUrSzHojrNmJPAXsGnxatqGU0f624C88Ms+WeNmgLUXIngX9rgAht0
XEeseKMhY0Ul08UjIbTk2aJmramR437Kgc1LB/yEuKbGknXPT41XmtI6Ebhy5FOT
LsKLSpZKhf7b7frjV+DQ66bxd2cI6zSfjmgZcnt/tmW/rfSMBhs/JLUZE6GoinZT
TW1vf2Y/GRGzSHpk3gPgF0Ca5EmPQDIzA/fSAebrAIx4j11bxieMaeZteFYBbcsz
LJgnkWC+dkF/HF/k9VkBlt8xBk/j96lb+UTmA4eeqxkbaKThnFKKszhD43lX8u0O
HS6FsTM3trWYt9ZtSWkJD/P4idhI6Iivy1wUo8is2FfanSDOobaB+c8c8ae7qDNC
ZyxT5h7Eu8cYsHZNgdo+o94zZQ/HCA8piLHI+l1W17FJjKV93RQT593OTP67Ca59
KGmQFfrKAZV3ummz/3SFew9e5/R5OefrmDWfhUUkNA5NKaKa08Z6Jf/ZGpHPdmqu
lS0uDZZNyXy5cJv8a98DR+9L5vTLhqgRky5YGrdObnUN/nUDLBKuzCT8zJVkgaeT
5hxdxTZS8z33NYt6L6/rcPMfEpACwLCciTeeogbDub9TP/Ur7J3GC2RYso5L2o2M
9d7y4TH0KLh1kCwBYBhl1AaXoL6+2WlsF6SUk7AUMxLzwC5+su2YKSNu1yAzlx35
tCjAvUzkuFvv9JNvdK6h0lgw8LAuBbqkIQQSad2WoVYMawJRDL+CK8rz6wwUV8/s
Nyk/dJgj+bPfsLAByUEZVEJYOsd9wMzAcMkRbsP+0fDKnWlVAu6Exb0h1M2ExAYH
0soTIvjWsxF5W7zm6jKBVySDkSg6HjSOFG/Ls+Sov6Rs4NAxpiV+5Pj54dLM6ClK
9LcZicj/1uyXdHR+iQDDZ4l8NO60P3zecOgOxgc8J6nDzOEhuskxvvRzmmeZ1ora
CYO61dfaTPZ8y4PrOyA7yK52mZDiSaG6BGEFKwZnDS8EQ0Bc7HNx1Wy8QzbhRduK
Dkos0SIVdE3Dtqc+HR/w5RyZv8mVTdM4OBAmT/AQi7i9t5xjyJAjnr3qO/+Oq80e
8uLoOjz90OX9ATvo4xXnmvVS1fu+f+7wCqljNYSJgdjYUiTRyM6UwKpcQrciXuwG
km2NQz6oKG+5QLWgtfrAW76TYsB9o43V+7g7MKBpqMYqRCg3XqTarMGvBdR01fzJ
ge5JzvnVHYWOOkUkXHPXZmXomy91t/u6Tz0pj9X2E2d2C9hVOvKT2w0PeojjVIyU
/iLbR+Xg0ifpbBFqKCjwBzeXf81/9A0NlAGc6mxZMenkm8xkeuncyppwCs91p/LM
oqD6MccNeoKD0XDxloHYpAo1nkqY1zkv2AVcBP3NiOe7Voy+iUniYr7IBoP/aMXz
zQgfGXbV4Xzp2P9lP+GTdjbzhDhiaqBolAvJxWd4vlaq4oJyko9oTsqFBdWXqc0J
KdecW7YSLpKnrueYCkmiGCinEEVcnsfo8kg6AKqVKrekpHiKdXLCPtTqABYT3BgV
5Viv7q6/AyyQ9BRKZaeQ9BmF7zUv+vj42RuWcLMShUu5Q4vMXeomgLmqSF7XmL9W
ikYDV46c4hGNoI4HbRgT5VKEe+KcbSlwk0uEX7n4FDMCHCBqZSi+RtY2v2aRtrgl
qzaKwC5My8BKpbbFfcXDtDPGsmpr/MasjAcp3gNpH8LGymkicbfMk4+T6Gkaggaz
FktpSD/0DUAZj7LdVs568eDoLCTnZbVgA4VvLTM1ExsTd1t6oG3/B0LIVAVo/f8F
90Aep6+U3DCQdET+2tv9IoimyLeCudIOB9BPDmyu/GaXaVbN69XBRqfZeyNiBAl/
fEP1taiBT6NkvZnPN98G2AOpvWOHgODc0kVA1xnprzxE1MtyAyCI5hV4POvbqM6H
Q44FB4jq8l2iLymiWWDkyCoPa+/GT3IOS9aqxSBjL1KcxID6cWfeyBKIN7OPJoiL
uW8g7M7yn0i7HHUoLLjtuRE8E4iv5r7IepfGMjq59I7CsfiHfA+ej1DbLLjyaqkt
SL8nw9lQGAoTplqP46cHTMCvekVSPn6yhxGIeZIFp78R0OlGWAT5eArbWoT3socj
VIOnb03pjvBNRsYsUO8W3kBKcwf9q2C8IUDMYxiW4EBvt8ZxJmYRjDnBmr/nw8ha
ZgW7g6qZROGpqjRdYFoFXrwLXN31pKL6OM/TtlUWY7mit5eHYXbrSvcYB1Rp4h1o
L1oy/6kK/GQdLrWHBl5jI4qbeOaR15H911m1J7LzggQG1+cqE2vTXiMhpaYo6azM
3KModoUuHbtAlRbB0+ThQpCkL8G/AH5lyn/cOTsHPVDdLq8hX+ULNTWZf2eHjzvI
CjFyPOgSIJzThtHphc4+q+BDuTjIxBLa2RAxNLFENnl5mJebQU27E8tGnaOPipPs
8cR4wJpfUIHqxgzeaZ6NPJNnIoE97AR8MyfUgbFM++yVUFg8pvvwUaYrweJlm0iz
Gym73zvMHtKrvc0EuDNi51gQwsC3ctJAdVMby/XTbMniaqkVuvWTYAeG3fh3OH8S
`pragma protect end_protected
