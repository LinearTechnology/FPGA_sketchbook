// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kxND2FIQeYhwJLLjYS8G8ETTHayNRdfMc+HbYCIlnV49Cq8iVzoVpp/mOzLxhCZC
Q0y+KtK+umOEFbp9o9Nc/RMK/TEi7eS8X72iJunG1pOYw1kmQ4BJJyvgMskoZKwt
CsqWyHnr2hgYvWjMp0qZxVYgHzPzxLeQU81OFLXELx0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 103600)
2fwWFD91rbc8VcY+snhOlgwxDsXJVhlVRNiStfc2ezraQqBHIRRo3xEJYLL3mHYe
F9OoGYiBJuvaOnoavzkGGi3c9VkhABBlDlPk1sQGXO7PwDEn3pWfrM2LQtSPAUkb
f9iBv9pTViqPbx1ozgqsE1sNrsmi4XVsVSvfAwq3RnuDpV/djNlvjiRj0zD3typv
xpHevZthH6JOkmOVdr8eFti1miwKMqXysxWI6JDv33fYwjP3tpU821HaPOPyT6RU
S4Go2uz8KpqsfT32IbmD+HLAGRYSwbonCQYU9iSd7SjQSmgcvzHnpGsQQvyx9RAn
fdKNKBbsPhBNMHy7FLWs7TifqC5Ki+SDPyf67G5u3zpJB9TvyU2pw8m3TrIZQd82
rW5PjFu4kssFsx+iPa4AXosP8cQGHOcTNrc49S/e+7nV+2/+UsA1nSwmJQtCXDQq
acAys35wZ4dDhSjSqS4Xe5G7p8jEMjVZEcPskgwKrf6u25wnbMaa/E+By6ens0gq
nSAiNbT7lNmr9txoYnXNnppiMdNR7LAMDYuLYSkXnPk1eNUacmdAfyp7b9iKg3BG
j66dAeWBLkAX+7m3vouxaKgTiuKIA3672SYowA7oQ9WMOVRtjxURDprm1bALrThM
fd8s6nDXOJ3MrxYHfRtrU5/r7RNXkM6l00UaqFEAFYr7EWdgwjz5LsCKTzB6+2gU
0mV6rs2hQhM348RPCQZ1YDjfi4/u/biTgP0aUAnZ91CtPUNeUURE64wwKp3BlGyt
uRER3KrnmEM2eOFZjMDTVX9Yla3bXvFrWIuQHXj2169fX55PBg68O1ab59bCVXGt
BC5smA3NJIF1CB4nsWSklQT8TXeCmz143M5gnBhShBHBt8ABJlRq0fj6kt5puWSU
1KO+vK3C77BqUleu5u8zsawA3cnoeGZqdK4Bs1GFHeCYrhNi2pVKFs9vqiSDQtjS
nh0yy94oncFVcYU4HJt0AdNOeIVi7qqMtF1rNZexbbJtM2PQPEjZY6CKKbIHOvIA
7Rbdtw/dZyjLtjwCzkUFooFNVjLDinOMzshskKU352OvgLMfqRBqqNx7E4XK818m
1uxUQ/7IK2Pv5f5AOzmS5j/9b8ky0YDFrsZtchwxgV4m40GIrQLJeWVhiiR6Qqv3
3rNbLHjGR+2f6PYoeBpy/V1vWoXW1QtIQya6QOjCQdHFw/8RFcl/qKMSeJx/+mAG
P0JocDhhL3PrSEex7K0rUL2K9Xl5LTIKnX06/pJNvs6Tkz8eMNchuOgkAlRTzuEW
X7FPPJNO10qVaSLnyQmsOikK+JgvJN41qnn6BA8zUK+19CMI/Y24O42d1vgwbCRw
2CkV2NgGvEjtAmL4HAKNA35oEfJvtP5UGmRogFUw5EaU8/ES0IZjTDVcR3sXvpke
M+/lVNpu+9ORqV1wkQwCK4LaIyqB/zf7YIFzhAdvAajaCoM1QaQp4HQ2WqZ8cai+
MBHjcWkfHvLFF0t5VcxuFY17qszNei+0yIBhZHTMia5gk3g6y//mAKpgT74PZ8Rp
JJTbBPZOOg59LkPXPeX0PC0CMDxzBjTdazeUFMsJiy/enctBVMWMNuUd2dnf3Db/
ZGMs6wT7JG3y8OXLymc61PvA1P+xYCufm3gAYYtfua9JlNp3vjs0eyki8u0zThKq
avu6mDLhBXXshzl+Sgbpp4zFE49+Td6lkMmKwio+geA7EdsEfNexkqRd/vjr7zBb
LT5jYYXqI5lmwqPMunp1dN+/ClnqKEQ18/7u1krj/W+woJ6cfH4JA+xvj/w2jzg0
VKJEgLnea3yH7Detk7qhU52tOVuewvAPAvSZ4iwMkwj2VuDIIW6q8BxOWnA+xcoT
+3ZGOgug+jAiKG1llxVT3p8dSCMFYuoQQfPo7uTkXbosEPLvIQui0wdU3KJuPoVx
ep3XPUjCkbh0jfbYo010WN2sGdCFp7hpMHIoNzX3+ISDqgKWzbm2yt4cbLsmP9Ql
II7/842JNtGX9FTOhv5iONlX7TF5iLPl6pB56B/Rxx9v6E8kEqwhG//Vbo6a+E9M
9+AdNooACzogWp7mlUBmcRRvvq/1H7rnexrldD9MS9oTilsspAHVAXqC+YYMWGEr
/lgI0/W2a1/ouxC1YZhjLanlgVupm1AJ8QTFSDOyvNFWW7pESQ5bbLD6X5n44Uh+
xJmvH9OQROSqAm3S419FKTGwBO5+T+OASsnYKZgzC0e0FxcUmGrtUJBRy4r3bV+G
zeJhUdRBZicW8Z7Ql+nurw477kYbQ9Tkg0PUzZd4jN3LY71rDAj2ap2JQ3/va6Qx
uMXOUVVmJAFoVcRLaEEaiSGrSUL8VMPOFDDUwNszGu08/vnboJMcs59Gh+2BsH3e
GvCLtt+sAt/bEMegjvxPX3oFMXX3lfx9JsePH3sLLHOkArVIixr2ea3I7PFAV/ix
Ezd24+U58M15/dG/ozmNYW5uqhmJpZxk6LQUW9CGUkJj+xe/a9fkw8MIIspJBz8u
hx7l9FwPJu0uJSbtQR8E6QeHyvFOQ0sUigMBSVfcGos6j8Y29byjITOqW9sQs3Ts
kO9AlMTaYkQXyvNJ+qaglSi6jCzfYMMtg1YMPCIlej72AN9D//L+N37xt8Es9ILm
2gyIWACHrh6qiIXx9gC9CPvGQsR+EEkDBR7jHT0T1IIw1ADTvqobzeE+K4jN+ZRL
v7GZ62Gv/nUgYAM40s+WGsPIOZPeJR+aHZOkyvVjaeMrdmoHe4/IIywvIK9yzUAg
1KcOCJ5C+1TlqATT4doRuPl5iG4lweTkxBFnHZ4l3Q8LzsP3Hx6NxwzjYxIukFnm
jz9DUTLP+tv0nZehXdBUGrE/6gRp3+1f4Wiq2PfxmdDO87CAoMWrCO94m9f0ZmdX
POeOywHIuRz/JZl0vGGhVJuFEa+RndRHERlG5pltpX4YaAkAEFnuq+WYmSjH1oX4
k9eUPAOlpKHjdZVVcegnZSI1JNvcEUD0sDLtUJozlc8ut9l75d+zLdmzAmhHpIvP
eEFO3je/n/CCW/f5CewkGlE9on4G6bkY/IM14uZoYoCTMkAAOnrdPb9UUt6CchiW
5nUyUGw9gAIKV4V3TLEG+fJnLaHIOQEIjWcP/+Lmtqc7AVu/8XoeyxRx/UFVK+Mk
TH6tJFfrhewNqRinSADgg8BTJNIFnomYgB0hTzPlXog2cooUcWDlp/lROajcZgHH
zFLO8p2HlpTMzIzMRcoPtctZcfNz2ddk+cpHQYM310IjoOdKSlDlC/psrldKLhmt
XjKeS1niGPIeY3UdwZbeH9/exjXtrUvtk4OZH+CSdg0PQzxqxV4giGVT+hMtwkhs
0uxJQpgVBjFoW1v0xGGlBGo5waKt5bVl7C2vJN4WmcrDctYfNEwkNLZW5C15JQHt
wHOpvwQ6MsjHtP1X5lBwSixxibwJVAFV3JESl0mA9GNUPgMfCQehqhqtOKG1DoA6
ANzTe4XHS3hfcRTSaJe8CrdTpW1B4ZbJ2TJnX8gVqcpTuSUMclCLrUkUoTfsZhwI
udNMNym1CJLm2fBSGdSEDYbhTEUxuf0V+YHkKCanZ/HlH4UrgUnQ8zKvJuO87rXu
HK6NTn3iZ6DClctDQA1HVRC3TknuCsphrCETpSGtFafxIQlD4Wf07o8RLGPtiDEa
x8cCwr6NfdDW0VRZoKz5H9s7xHK52Gv57rJ0FmFzIHyhOWhcGSVlhDhRRJSAVELP
yfiZLp9U5WVENfUzd5J1N8bfSYFbTRDWJ+PUQeFlAki7Gq7ISH9BkU5YefdFuUXb
w7hMTMdAfvGB15+gFDspigdjcydHR6E2uxmSULur/JmZo0DDffnXTNZCzX+6TDqs
2xdTvQJoxDIYqHfG9iZ/WrmTx4EUY59waZsAKPrqT5HQDkuRRXdynFavvELXP+33
9GYu8hX1pEJKHLGfFttZUTTtDlWtx+stSziSw5+MgOdJ4XlMzF7vLzPrLix1r5vA
5oM53JM8NzyvL6JxdRRssIcVDhy8B3T4PKJtvHV9ANbDFowHGIuHE1EUv9Md+BQM
stC2x7tgg3dl5QjeQZzNtO5jLP2oU6GhnVmkXcMgoCuxUxHH5EyyPMXDOHj+wkY4
BfmGXLKWyOfAMXJTNG0TXa4mY4UMMp5s7fxe3gBy/Or7EJrga74d2lWqJK1m2XkQ
4XJqHUR8Rdortem4U1h0BHIwEK+dL4T4aHPNmz1ne5Q8g12xaGjkdb6CIfceHoII
ZSKQUeI1p56HToQLB3tzWnGCEekkBH8pfGol11pWRwR0En58oRSIrvmI1sLiibm7
vyaSRE0J9Hn5mzwGEJccP5PQJPizVTZ6i9ytY1wMNTf3WuPmPjSf3I2K7HtXujWq
ITZGnCjxkzfadSwrgtB4Nlxqsmj9YLHM/AI+aIqMJ7exhJTeK/JWxUY4j/RCQ8nW
O1OwuA+wuIE5LP7PXIu7TvtaElnDi+rmy0L4TJXZMD2T3ehaNVF7MYku8NSmyMXE
4NERd/gTitux/ODq8rGI7y38kNT1lmc2ezr1m7VMOfkcak/6mfRk6/lHipfnSNLx
uCNamHxgFI8DWZlJ77G1kFAvotDMFt64XGofw4fRDD38LoB7vH8QKD3zADX7RfFY
fJZTQIF9kQpz3O4+Uy+BTQVJsqRW4PDwWRKZlvhitjKKDlusagrYwnjlxMwMlPwc
TamyNiBdXl4pumicG01rpVje0uCxP+BZ/+lEaj/eyNjfAle4Jsvh0dHGKf7+jP20
xX+p3mw5nkIFtqVJGwlBb89wO8BMkQ3QbH5wLPxzLg0wIZfDy4/FRwfdT4IYCEHo
FpLh+lZfpDywHHFgFKQ13n+J/Tb7oRMU0Dkm9E9onRL42v+PgO51qw+Q7WIwj0i1
sDcR3ViuA2elwexDBbAURnQ/KM6DnvPFRQsW4DujQ5um4gQ0Faygu/K2rYnvuQEs
jkmacF0ML4Tgqwl7s5a/zosal1KNnWlQcpXYPFxnG8n8nJ9ZFyDkOhq+6JLa/px7
LgtVQx3KoQm/mFvf868aXJXzOM/oXOQ+4HcPMzhxB3KqOBq9BMdAwxp4+1bwFQgP
aIKX+nGzZJlbI7td4FUxGPLU+f9r3tzDSBPOc4wlw8s/BHFCdzXM+SZmglGhn9HI
kqQDMekuRxMLM/RpdLotkGniKpoSM4TAazXsXmBZGZnx7gkbb1Yrvm1BzSveHe35
opD15XMs0I1dA9y3EO+C7G6JH7ZWk+v5XxL5Hl2u1oH84HdDbN0k/eJaLINqk8C5
xC8qbRA2FQz18dnsUpjlUrYwqDrdfIxmnGlK5gVY+IdBrLjTljCX6r5yja/4g4W3
Nbk+NrlJcywvqI7bCnS41mg9JnxeMcwaJoFU3DxM8oqzpqzFsdFknCNZkiTBFS+z
odRi4naII9et05MMuXnlhPb1JiueSh4o4UBSwL0lwWVle9QGguDN4CAtWbgAvGKB
pUt7pttohtKHRlKdFZjz5rKvC0pUsAs2ZPD4qnfR4SFegDG6S+v5FyoWPvwZj4gf
4AMk6t0uYBGWteTC0z3TZ5ctaOpe6mLXfiRx9pA90XyDuoKQOBI8LWW96vRUWFOk
i8mnUdRV/PUa9GDEzDqNjmyVIwyt6PuI5G7vIreXIzbPIviN0Of/inIgvDT82zbS
/44wlujmkzYkdjb0f6UfMkh7gFaeeeQGxjNNbWtGymCriTSj+1iJldo9sEKB0PGY
ZYH13T0oQU7Vg7QXBq62te+oC7FB87XS0WTI6aw7dVK3XPAyMe2t9sVSA7e5H98A
tErjFOIDmGhzyRDEegT8w/I/tRp0SAKEp8Q4anFqLG+v2DcSUlD8tAgyluSS5fFk
11Tvp/tWWmailErFExiGrPNND6wnjZCJ3T/J01a6YZq3ZtIjNUJiNsd2SlqSruHC
8IFIcdamxNDt7qpqKpzEv09wFeR4kiBabTeNDDdfiCsxzGn02WU6fdaubLNM4oex
xcMVjjqtFwSto6bxuHKGJYUbD3hTXD0YVcu+slXv/B69Ed0erAEaszslFt5uuKLl
Tlfd742qWYjSsdR4vdzpFeX3+VtPj/Y+9ko0QOIWh0IBkvtE2WeaidsV4tMabAkf
B05cM06wOqb2/vTGPIhgdxBR2/kOm4v0+ijoXJ+RgBeabffCtBFRuAG+NL4kMHWT
9kvHojFVI24qunDO6KEdo4cVs4qI2r1FjR9mR5IihGVOPbRfMUk5pZM5KZC6Mbga
g3pCF0if3x2DF5BmNRWm2foCALftsZCCBV3unNPodhk7NbuCMnRj+2mhmN+X2FnB
P0yc6sEahuO3vWDAOja/7ex4zpVLrBYkwnsx2rpw6zdNUUhXesi96A8xnjH8ho9O
Wt/fqBkJW9nNpETcNUq/KafijOEpbZpkKjfYncHQshhEh6PAtL6u7+C6y9rtdP52
6XdjlTQIjYvd8tfDUHzI92A8LUr8fwkzXsIZ8mj1nDb/eOxLbT8VDp3r7+vFqdAJ
JDftWnaFNowwezwqil0DIGVl1akE9Ci5680C85WvQVRPYy3/ToC4L65lHz8fZHoi
a+Gji1sY5vkXNaCrLx1HMhdIVpOuFlfIz4McoR4bWzEJ5fXrQl41pAjXrdTSFLMf
/V9ecT/ufopTJqj/mn10vFg01PII+8rT+ln7HxRRoNHY7mju6fIwnwpFqz2CaL6J
IUzU6T5gWVpL/T3U/uRm1wMVsrS/u+fJWsFy2PULxAlA5W9gw60PzlIGsW1S7Z3v
q67PdEdmqHFu8nxNf9/VG98oVVKgdDCfVPEVA5S0tYLMUrtVCXEARtuaCv50wDl7
oaR6RicwyNSp5OC6rEvyT9vP8QggRFwSsWY19tqbj8luzqnjTRW9NfdTU4EThIrs
4RlyfiTUo67u2Mv1e+nOb+Z/wfDJsYhoAq6H7+zqoxgP302SF5K78AdIagBHRIc7
hNoVTK/16a1EzHWTn0dihseJdoSHs31mQsiOXSRH5BI4Kz4Ax6st+BXYX8HfAyRq
PyZ45WSJ1VaEoa3vTgAIJOpLzYOg92hsDaMEnu0PJuJPSqpjn5jRz3gx/ww/3ZjH
Ey66o/SqWfN/CInMYx6LVB22+QyclnTqGGk0nPrnZ/q387vWY2/egjGaHiEgSall
l/lGgKOGGbEZAOsTqRF4NE+7YjPuNfL1lp7v+dbAgGmAOo0Y6hKDrBd8IEHTkDZe
nO5JZz0LGHdBmElvmVKBGT0lCXoaLw3pgnEhsJz1innrNlN4UEcbXAiesLMp0XmR
kYpjLUcnR1KQDEdQOeiNUfC3FTRNo8MKSY/7uMUK22hF81aleQ+r4UQzjObn2nSa
z0arqWt37z6WVSHsdoA+4YsppOV52UtiT0DPN+1q+sg93lB/e5NvH9MiNVZhpCPC
jA18JN3r/yy+cu14TjWBtMNYj4VQvUBzxXM18paQed0s4FsNcJ6CnDbyqJ2T5MUT
EqorVtTzdm5kUcWoeNVZSptZivMbSZdciKkzNx1GkMlbsuatpXM/ueh/H7ZtBsjX
YS78XeDKLPAiQnRvEB3nYWjXgQHP3Yor/Ps6DSweyutX5EmU5KuywT9yKFNfpKzo
9ghLUTQ0pSkvxjXHZzHZlcxmKn/OSMHNz2ehSpj/S9HWNmvJaY9u6mhSxKCRQz+r
yUKKqWw1OWvBX7tu2WFHfn2nZCBWUo3mBxXtXZl0GN2uNp857DVjMb+yZAXyj4UE
/ss4wTfoXYEMUhFAwA8zA38MG626fo9laC1qnuMKnXxaOV4VF9Hw8f+vsSEDPkn+
+TIl9vBe3ZgiCQySVfi+jwkRprgoOF4l+LpiG8fKuwlMJJeWbxbjQUPUdS46J+om
+3ToNmpiWjyY13rk9wTokfHiTW215zRelEyxZlhTYYQmAhVrDmJ+vlRF16ile2Ag
/UoA1bT0msNmaT6LeATyfgV0rZAcE9Zohs4jp2HpvU+fkR3JXotv9AWt+vepLsJf
p1Oykm37Pgimz8u40pCpOM3FfVkH4UTpiP7LOaWhRp8TWyiU/24zd/Mjm+Vt77iB
DN7VcJX7zAml2bDK8YeyDHIujwFv6rgv8l/bS00nYUOQYO7xFxatZ3mEXpgdbqZV
an9hjryE7skFgBX8E/2VUcQZq0dMr8VHlGkWA4KXishncQL5hg3t3NGmAiFykDgc
iaoUsuQD6cyEGVCXF7GQtGD2hN1CixD/hkdUcBXt9B8n/dS1TXn0AxdShs7K7d6s
Jzk+KWfq3Sz89DHxOU6nEdwizuiUEaoVUGYXTnYoOxdO6d7mFSCjdHXsNebjUdBx
3YEsS4zeIVLS7Z36nu8VltsF5FrDn3pXJWMHclqHWT+TuUMJA+VogSotJjGrUusa
Of4yH782bBB0S5A7DwimVjYgBGU30GtKfaSfOH3MRRsnO4a9WL/ol6otbubiEm3b
F5ZcgJGQtrd0mLcA6eF2WLlNymkxplFv9RJQL9oTKZ+4yrsYjh4BVptxuoGfkoEU
CQjH7OQ3COHbmaSKrdj9xaCqYJKf0P3M1l3tpQZSAcnVeQRWxLX2zqnG3j8GBbKX
+SFazXeNGhbpfTkc0iVLzjJ/Zy/4efQAqWUdpUKDh4MPzWhzy4jgfgwgAr/Ey7cP
l3pPuN8zhJJ5aND1j4z8+3t2qkWYMJ4EEJCUEJRoHIwreUPsqn5udwsx4B80C97f
8RaH8d/T9d2YvUUBwAS4UuBhm8oWg+VZKznWtQJ+kIbEU2JruiFQMPQUf2HYoPpr
sQVz1O80C4X5qRdchzsgtXOEDc8257vl8lF70padareaxyfy1erlBAvH6ouJ2nUO
Y1cH7gHztGj+jhoUPizqd00I3T16iKbPQQ/P89jechP6V4tX8xu2MlTaQ3vRNY1f
Y7SVcZvNKmIrYyfDq7r8ZVJFOk4tXMF/HAedY9QZoU/8tKxqw/QiHJwx5BYBZy3n
T+Io0X8xGhEH3H+NmxhXb/pGhL4d6COATH2ttX06thSd14DNT/YtdhcTeEEJwTSE
CA46kmjxnMWEyGv+dIMynDP3a4dy/t1CUYFuYQtbpTlwxI55KkNGA/GkHqzJQQ1C
PcSxQA5YZllDZzGRNmNa9niyYthz9MJxGybviWUfVXzPZ+y2vmlLtR7kq41FM/jx
b0gjQia07NAUlQKpUOnl63f1KNvLyr9OBvwXMQZIFuoadhtBCtCUfVFGE2VR5zdY
62zUmlIFlk6FXWJpXgsSFGL4REjQXnTyZaO4HYo/AcrWxO8BMS9cmOXqQRvyePYr
H4SH4lYQBgbrlmJgz4s7aEo2JR1YsRtLkkwL/kmYIpJZhBkjzn72rejtNrb4LCoL
t0VMx15nT7UP65TJG+8ow7gIJNPuDXz7uuiCrgX2jhnCcz7n9aaiekYnCFnEKoGE
B6voPPHf/p/R6LBG/1++Ur8MPg091BRvIRH8WaNlyAO6Nshu8dOp+G9tmObGPsC2
oS5NH9ZbTLDsRKjBr5IqrBk7CjADMOZ2+wLQVmCGKH9Mqwjc/vIUluUaMfo/z8cv
6hRd0rQfHPKxOgi7B/dLLmSkMPcgprwc8O6+5cS0+sMfLMc3JuHd0F3D2UGbEsT0
YopdvzGcpJ10SeIP6CjbjQT6iIj8jw0XTLXwYeTcKF96hiEC+fErvUuWy3p13qtZ
urxtK27FMmNeHPivcXy1pV0nQcIifTEH5JpBhKkWUOjM+Yc7x8naw6u6VJ+5hsvA
tLXbCb6UUkOySMTYw5CUwVRUXajtedwso/1CQ/+Y9BM1J8yw29YCDp7nNGSlL8GL
qVvdKDJuPeIubp+rCJYv+kkT/p9d7OSiC0j/viSKA1BwGJ37sccmwuobiAYgwfn2
oYwbbguSFfiQaZbYnYtmRGvCp1/9OWYeyBmmCVb8UcUuyd/kIKyK/8AElPvx14IF
KQpg7Ap3juFxbvWJ+Rk1HgRPPiJxhTBkc3e6GnuDwaaZY2DRZ58tlRKY7eLMd5Qg
PkKznhzH/w8q9nTGC/7xtkQn/qeVRHvx1Y3VusLDnw6sjUX3AvCzwSoxWKH3+rkP
+TwhtEbiPLEDspuz5Kz/axF4KyJSxUjZQpopstIHHJDgYdJmFEBWQe+SOatC7pe3
/x0fxIGb9DcXSkrXpBi0QP6Oyx0AE1z82m9fgks3PQCiIngkQPECZFX06msF8vKh
wkzPJbmXbIlLeZfqLkP/T7SI/uHxDxSmWnuXYp5ZMtkiSfTejJLFz8ODTKjwD870
EJ4/K8pZomvQQxZC0wCBBZvzBW2nXKHqyAf+OQM8azw3tO82mkVTa0Nl0BHEKNFN
3hPNKlThu/s26SEb32mAxhjNNVw4Ekgau81j1ZoB9xDczDJb23zgGIu9SO7/NQ39
GQoBarLdM17lYLivH8wki4tqnK42NQJRRRWM68MdgElevm2x3EsVJYCUp9j4R/XB
j88WRXAxz9pTl4V+5vZ5zxXYUJV22b+wjDFWNCNyuR+Tcnk9XhnrLTPlYYkeLCQ9
ZkEMKQg+HwpLyTaiGeG+mLiIGwLYtnzGzIHBsrW92N8rv9asLQUY94T5eoTiVxl3
pwNsrlSdwS68ZYjoR1zrpmBzGu9eZzG06WYqb8ikW3r65MPGW3bwBVMIvWD9oHuR
eoHnjtNx5i4eOYxlCFGtguZ6hc2WWJNlW6h05YMcsh+Lbn311tL8+Q2eFLDSFWrB
3SdDPKJEXKeY6g/AvY3A+cYfvPXG70t2EcfS5TGDYxa8Bk0jMMFJwhy3KMjffbrp
kI74kJlNK49CtgVMCp2gTgGB17helm1juYEqaVecKilE4jbUaPyccmeeWgmHKOAO
7qbY0KX78eVKGtDmQD6bgbSJ9DRxgDQjSR/LBY04Biso8oBpMeRXlTkLLVYgQyTP
SvpA8PE4FHubESY6dWC8iXJywJAKnDraTMg9Hk0YRwOImL7x1J1RyNYeEVV4EQOn
fwYe7bPLjg2I6hzPyfQmwgyUk4cMCfPKNnxAaHmKHtOyEbKJyjLjYJ40raamA8AA
JILOSsgdJVVap2KIyzh8V8lfyX8O8AkKe/mFd2xkBViKI7J94hjytmHAtFuKVdQt
zcy3EfmY+b3MwoKUEq0k4cpmUqlh0CYs4Jqio9V0mEze2vQpNUlI7AQuiC3m9o6/
u0WDepCdgpL5r2nlgUao2bM6BkLRqCwkoY9qNL5cN8U0QFS9GQsugmq9qxLrOL0z
4m2F36qQROurYRwtFQ6NFRrmZCNDoTyGNrknuQrl7JkVGLNiHeV26C+l+4xgIfRV
9JTxPlCqW24/UHfEYX5O7bAWqbrKFZVO/puBTkdYF930roq7NEstRewjoYB6UfJN
mdCcQ/7LZ2IJ+Ynw4UiMX9slTDauwCDuRQDA+YHV651LScKqCurg5vlPzT97S2Q9
c3bUSbItU8XhrHdyWDNnN9/KArLy8d5my6aEZ0Mntui1XcYL/sGS3zzGV1E3kZ+R
4l0fFJxkumG76Wns6TPf9bWWx3ro4XBA9WgPk4eIGL3qryTLMJz3f8VamtoHqFZB
9ZS29D6S0ZQ/HCxSHT9ZGV9yyAeeEru0U2ET1Ld+a/TzQYI72pJq/18y80j564JH
ETkArkQBMHK1dCPNb61LJVNNZEeB+JGZrdZFrIrKXhmnpkUx7e258sBMdqI30znY
KRDzOsjBVNSHROtV/Mdw73n1LL862TWvQf1Gxl2ae9RuehLQ/O7Ooxb+M/qdv3oB
77t4gLzbDNQTvvZgjICwi83Uthu4mAcTe0NinJdcgm4qa9S7LSWVgDOVoYHKQr/T
HRIIO3pWHGaLpHH6n4pgYmA0ws8W7kUMN3KejmyMY/KuUX3DpRihNhi+puQ8oziz
+dde7w1PWggErUAcRGQkf+lgye9lNY13Yg2o2wTvgpkIkRtVobWNTjTvz5bIouW8
aY7v/8kA+Nc8LQJ8FgJBC5Al6+1wicXFV6xs3NmWyklo0rGpKoZJGUtqtFtyRtMq
8YvDNGR3VzB3A+hXE4svNmCqyFiTd7QZzvLIzHpx5yVWtbuFRf6yEcX9bCbHuv5a
UBQPjEqLfAtrvtry1SBYx43u28MUHVuA8tFA/4BlSDPUbEafCFWun3isD4tE0+HB
3Fh7obqQXxJf3ExcwaZxST3ibcfB0W2bPCKbu3DlMAUw+RHblpV+awUo0A0tEYD7
HHO0g+s1I8eq8REBycNA52XpSGbIpWEUZAfB2r/B2O3OOnXJ/CO8Mfnaa9x6aoze
R9ZUyTT36I41QYYbaqXTKKZWL3e8KVHejlA8pluC97AMdJM8wjbTWHW+SoIXkv4Z
Ix3Ehs2qtvg3STtmgMxa13W8wE9xay5VuxlyfTI5PmnacSCANyJZ9+jq2tRCG8PF
xYo5x3NfLMDjL93QOcdud8gpCqLncjjY3H4NMNsqEkAkkat5V8NKyqtcmGS9/gYk
2BhOkpGzxOvE9VbTc8aPnBK9GTfCTbopMeR0WF0CKAYUCLPmQDyHKwdlnuKBAwTC
9dU2DXvdwEbf2A5k0BQk+r5UuP8+80cjKQ/p9K9OPPmwjO95NmJCuV8YPcp3879N
694cRqrs1rq3pDaQa8+eSCaGWYo3TZDyn9emcHbJz3X37YyB8KkPUVewO5wNkuME
hVtKQJQUDyLhpEMvp9R39aSpAegZSzNyX7Qdp4veyPaRL0PoG1qNsXa1LIfbGwlM
Rd/xpiYQzpBdnk4Uiig1y6uy306YXHLDF3k69PDRRPFjjewOSiAMwvvnnORJtOk/
pMHZfyNpMBCE0iMZaFyeHhNapGxPDhG/ZKLGUlRbFie9uYkhwO146y6W/A4NNRBH
OyOmevW0UVOugcGhyPImyYKxkVPWjwu9FdUut7td8a3Tjd8JjwESa3wwwi06Kpwz
GF0ZmwSwKHlpTuSG1Z0PWZmRbAd4iVA5sYux6IWRRTBrLis7wwxiVn4pEI0W/3r8
0xtTns6xd/4QQwqWPSEYoQuTsQqpBzvS9cIQopG47RzLE3xMTRQjBaeEVYQ5aHgT
fcCslXOxhIgIlZfW6RKxr2mjzn+gpyQn+LRqhwDhKYtKTiD3QST+8iqVFSS2wTS0
OhDhozTXfuq7coxQvydZsyLb9fspNN+6/6L3x3mULSIZ/ucV2WfgElNuaHJpIscU
my3n8YJhiAGuIx3xG5HAdLuA52/uBeOrdisAaWdc33kfmoYDhVIlwH9Hvr23fyQh
h8z2lGpOkFi/C8qK0QRn66XLbysVMYvM7cdGDLN7U62Q3RwxFbVkMOveQh7W3iY8
PHuDqff4S1MsN0r4tZUyvMmjFZaPj/nErDpzriFqrrSv+D4i5T7vGQ7v1rVpfaLW
Viq3+I2TYh5pRSlrTLavf4mK+2/sRVGc0ghYPhVHeZPQ799BRKawCTlxLxK1nO/M
UKMOzBDo8kr427eopL+ywap4X6WGmNh5IyulIEKFnccSgdmUymaHi46JUU3DArQm
AR79KBEDldRZnjDveiADRJ73ovJChBTs6IuhcyL8ggjH9/SQI9OHBdmKfEg59xo0
UM1fa8DYDBNHy5S0n6D/tPDlsDcnXX+UjFWLv8elYgZn7QCp0Y0AqfbP7Gqc1ucT
2kX1z+oTf8rBvIYrGpj50wE8WYoEvuKEdkRqsp0lidlk2uZ6rfAvqso7YVtokzKm
qPRle6LdaH2jb0Sj4YZ0jZbah5v3rwX8vSqxbSVs3qq3DcygGWcsKIJhypxXITOe
h/yxzHhN/YOPGQvmMPsNtDIbztbHC3nrf0QvnwLgpGnkJawznag8nYhZTjCL2C67
dYkfxtIrQq7xH1U1vWyCrFaQtq4a+PtTm+xemkNlTfwsMqKc2aHKb8mf5k7K2cfs
ISCwdyfnE5VfvqSHeK4679TkxbyjTg3Pz+hL03ackedTeR1S1FoF3rKFvKfGjNPv
7w5y8lbwyOMrmkIdCuYBWgVc/RhnK9ndK8UggVMYzDqVt6wiyCNs0C6jgAVjyrfr
1lKQpbAAv7fSVnYQ2AIxPtH6MfRVx0IC0RWbgid5IY/5qkTaI3pttao4+RhupGqs
p/stdpZgQik3FwIbEw0no/c1BXoo/PdKdP91+zYLzlw3/Fp2TSKKmlKxf02ZsYTA
8NBodtsxMoV44W0/4vjVyxxw4RgWXimouJovUkYh5Ry6r7gw9834IgK4QdGaIvRQ
6Zx8BsQGCP5+Hl4hBebq057wEDGw+1jHRCbczVNDImqSpwKr9cv5hOGOsywCRqgj
fmo/FTnNQscTSIUbMdtuB2CjWaq7TJSUtPj7y2keeir42Vz0PZ8JsrVYndFfu9hy
9WBxG3EZSGUu9wbxaSD//JH7r3ZakMG62EqsTRc1MuRFtq5qKGAriZ7yz+AzICbq
jFbn7GLID09UP9kS3xdnjWK4gKmn9I9TF4K2dwMs+7Grm9gAe25fR/MuDD+pMQOn
O7QePs9AjOvAVVCq0LhTfdQEsuJF0WB/xAITQMAHkn5bLJvAw0qnm6BuFAgqTGfQ
Rz8b0cin+xf7yEBmfc1AiqMRFGZJEN+cEZWOt5c/+XlPNYXPymN9wRgEiWuUyn+3
Qor3IjXTwEgnHM09YqjlM4xO7yTs6FSJT5sIkXeb7G3EIldx6Be8QPlx5jRH0UAd
3zcuIZ61z8325ISrFYoUjNogNJDKBdlf398c1X3SQHSX9G0vINndE8w3R4oibAZ4
W2PNe40d2mQRQv7F9eg1IZIQuW46h44AD4mLoKnCCmiJ7WnqxofiRdqoQLzx066k
7S4XEUnh8Z5leYWUohldAQTKnoJc06LubqoAB5ENTm97lgVFj11U1A58xir0AMLU
KPXPQBDziDe7M1CWk7nzGzB7Oj2CUTDHaEOM+G0yhCHeSfiVWDFTAbdsPzMCLH6n
P2xYGkPC8gLOHqSskafV9WlllNVohKs2Ng6riYjp757WXGncDYetJuqOppWkpr7Q
nixGRcQEC6K0j5Qu2L6fbOrxVRfeMTvssXEU0VzHHGRYuYCkgK4bfoHWWlx7OHQK
n1uZRAaKQ+Sz+7PFks+8E8J52ex8NOY+vBEzOUAyDJEJ8cZ4y2Bq5ErkXNOQJFWR
zeuOMDYB69imov8H3JBSRloa8ZLqVtdt+84pfHwCoLuLrjG8UFgoy2oofjUO0sEV
6E2RvMTRM5aOsg26KkKUnik4wanmaFRFojWAMyf+QjFQE96mMjiwjPwC6cB+yeNK
v0sUS2WC8jQrQi0mPoXN8mVVZXMecbdfayxK8TDV/ikRpiButPtCHEn6cEOIDZZP
RfC4ah+Vx6F9Lrj1Utkl+iFvCFtQ/buwz6ANuyM3hIN1xNKvpviSnYZ7revIGrnb
622247TKP6yfvdkRJf7uH7RrNFEzq+RVQoFU+L18oX3Srl55amJuKSEM9nzSqZ8U
6QfAtk68FSmxjtQzaQkMUeJs1wLO1GCkDQhXOS5rzruF23761N377EbMf93Efi0x
W5NNxJJmvhAUntviwu8FAGt/UK/xwencdJKlpo1ISbbFjaGDzIaOQHDNwJn5GMur
z+qvltbu1Keu5IULpUTjvScj3C+IjE2ELzzNkmXNEuTENmP8geHGo8MyhGYMBzQq
xw95L+++OMhE2JXyqjdxS9vdfqg2Q8h2vkJAbU83lseBX39qgirQ5BQ/W/smWoBE
upnVgHyTFaKSZcOnqHcoR0e4UfrDh7D1oUpYUOsFZlgyCV5MOeodbisHFEVcy2kD
JNJ/aGbjN7Ma4+b+zc0nkdtGw1tNH8GyEA+D5fGL4Sx4oSq3et4kyfRUN/2AqzFS
weSelXDxuUMuB80S6ZT/7XAqzDQ8efnjT/yYPPjWN3kLdVBEoDLSGdW757EMzmyn
6ceGLa1idCqt4vaBFQ7iSNfPfpKUKYStt1iIxdRwFH+c3S1GO+9oVf+lz2JvXv9p
WlbtgbpRR0/QqCZWvbRXEvF++JW30hR7mVk/tcL4fSH8tDyTFBIgeRFdQrdH1nyg
BT4FkYTJp1FDQPAMPv6wg3y33KxMJTabg5ETBHkD90i5qoKaO2TERvVIw78FArR+
a/xaixGzlRzg8s7sygS1GEuC46ANPNt+gaNlaZDbk4HoGlVsYs9eei0sgIXIjzGp
nmGa4sPf/mTYV+eNqrtvlemjkCw98G8wAoDht2+5lrojnsI16Q0OmJv5TmS2pa4a
G7sEoBNVi5WxNBLiQA+Li7xZJfLl74ahLtLXGeOlXITBc2CbR0m2dcwcMXOAjVQL
9WDqD4X7e4tu1TupXcwVzxYt8vVzuZcxcsMA3LZUOU00cp/syrXSVNvTX7AWJuu+
WTpdkj2B/4Yu1iRNJCgTubdXQ44Oln+H9ftdpErksRgumFRHU9WYtRzaDeVQrOZw
Z9nETOXejdgVeOkOllZofPvazPCBaIatsF4P5tT4ucsKoB2ahq9rhWhEzj0BqZih
qnAAGalFxYHUllQLUDlwrYw8EHRaykAR1Y1eGYNQ9R7ZLOSS3MbQiSQ22NXwF06L
cNGL1caAsXIKjzbqNBmnt7PHMmQftktbsMxW8MzAsq92wVnnDA1io14eiDvDBy92
rhuRdZjL3loArr+1graiGfbjmnfhV+MAudDTuqfOfcBS93FkmxK5z09jZ2ogch57
Xlv3zAL6/PNk6EOC0N7jXUZ9s+OpVjLcuoteo7ccfnidtaLNMbR8z1/Xwrb2pbln
UgrD4l/KqiErHrwj3EJLq9WaKYW4kZvGp52Zc64NY3WOCWnI5WlWfjNklN1KBpSE
Wb2sDUJuVYY2mk+PvlTIuKsJatWV6OnHIwW77v/D1+0JX/dcPqD9Q9LN4T99aPMr
kVTV7pas77cUwOdxbIn+FYsh1JVPW1tAD4cgSMVGuSiTqfutA2QwyR50hp2wpWw+
b2tyNgDn8KIy/EOXoTaikJI0Ox3/qdLZT79g2ALnVSaMDUaM3kZ1cIrWjykt3UcP
x+J0lcLyNxA6tdSsW/KOYNUhE7oZPJnkdWuSMpqoOcHB8hwgHCiuoK5nPOF36Mxr
nMn2sYq8mTF32EtHZblubaSsobLhpDS+KhlMgKrfGj/eb356MFvM3JWBBdjiGcs1
8zCwDIjiV+EGQzNmjNam1mV8uymrjKVCPSrblmLLCKjdCChZvo5x8jxCHHa986aI
GDq1jEGtqTFefxNj6U2Czf2lT0Dzo3LOaC0YsVz9nZ2OiT1temUcXZGzbCh920WM
Gu6bnCq3mq9BpC4Q9IYXGzZTOzqLpgdJwc7Yr7Mc5x3pvMATMIO/Z6wdqcR6rrzI
01d+izWbvQS0/VdJ7OYM3kJVbHWBI1f9TA1b0D7LCFD8EAXw/QT/YcKqu8DMayea
91Yy/9kURTwHIvW5X753P8mmr1nxEFgN1WJNQ8TnPEHlXYdnVYHWTNOLevEJZJFl
niDi/97DxFLpucl1SH0nld1Q2LVkMlwvjHNYTw/S/6I280ykkjG5Q9j3LAk7V9aK
1l+2fqsCOYQyh/rKyWhIgq8Ju6VOEXPOlkNeDLF/apS2aviU5bZ/vl8GaLR7zLbR
V0Ox1CiAbQ5si/ZYkYAeL1TRN2acjYxmOhLs3grAauzNxaXRLHGDubFXifuVjsO/
NROtSAESlOLLeTLWqYzcPEcbgzCD+6FEZrkpInVcoTeU5nEInDgr2yd/bx9oRS40
1csH2VGHf+ne3tmekgB8SZ73LIrKKrfQu9h1H0Vnj3KVODPrGM12PsEVHm6uybm1
IfAlHvBRfVyCD/hU5r+nkZ/uzVDx28ZMehgUf5BcYmz+YwHc0lJ1qtbj/t/nK787
XhZNR+x7kxCnPBgC3pyOYdgndSDFecY4l2wxNc+JPgNPWqFM8RDCla3wAm1+znQB
Uk6b42doa8JUkc51dgW32wGxVweUOp9Izv8cBZ4Ohxh07VM5tw7z1nndOuM+/gsH
9+BMRs/qc5cUcPofPGrHQLoLzhna2lNpLVMZc6uuvWy9/raPAL9EfxG1fLUZ1or0
pRCUctLMeBW5hVVCT9krhQgDjkPEhyDrXLD1jWaY0KlhvBxEKK3PKRVB4Ii9QE5j
8ol76fHnoU15bMhku0HK4V3hse8O1aHByOzRuaSWu/tyGkbAvs241VlWLJ9+JIFb
FOnzPCAw317ONSCQlqGuNyQqI/I6Ck8uwrXspH8nfq2KCeG/ZDpsuFWt3q8/GxNw
hpJ/LEYRXSi1am4UOIu5F9CB5w+c9dsaPsrj2oSwKQZOKubn2JfWaVXiefeL3wk2
GSvmHNx12lHU6tm+r25g44gnLoJwXZchDZtWyVpPtmgTM17icAlxNIuZjYcr2JcJ
rBzQSjD6TETIXrxKmG5wqH3MFcuB3KQ80rI7LqFnwwcRht7Fh2YaviaEuHf3Utoc
X4te6K8n170CdGpVI9D5DaQZwuBjluXm0/DnLi0qTRswY+42kgsT3eQu9+nGdNaZ
vWzVdfoACmuWYoK6dqsmb7kY3LJepM7hZ6MLl0Y+IUsbxwJ3qEb4femh1+PYp65w
Xp8YPQRxvlMMMKHGWZvsBxy7+8jwX5vZKygATtIV18gMtXL4dc5ZQj49wC9S9f48
8ORC/kY02YtTxJs536pmRUhG+TTIEp2oceXFbwKrPAAmOg5QOtBFl9O6hCPgQ8TC
N2Zz+h3OHSJCrn6HowQHrneUyHQ3sze248BB+cX6MsfyrqklvRr5VCqIXUpCLXuh
Ybdbke3ftrVVbfMueZZKVPsytDjAswdaK0tsf7vUNXlYBkOzRNNAI+GIUurrMKY1
EMqSosXCk0wjYeLgNL2ToH0ukjResK5GktCwj09mFPqqarpDibdUl5oulDhz7Agf
A6LKPC1LWQPQjbHQP2f0Ta2RLp0x1wUmw0deMlNcfKfasrypxU7AWzwIAvinnCFq
LwfStPd9L/5ztD4gOnthrEAsicbUApFIK81CP2lrBl8v3OB0QPIsmTE/SkkelSj/
04HlmnPrxIS06I+L2u+vUf126q15C5jcuhPROs3k9g1zvurnK2PmkH3TGzITngzu
rCJ3xF/RcgBL9lcujJs993xKgs4L2pQOESVJO2HiVwbWXQOw47UN+8HVgHEXBFgT
FribrnJtLJFw7zd951gvmlHcGWbB8T8lMQ/fpLeDTJTHnF/lwiXms4Vx7Iewng7k
nxzSGe6IYwAIIKIu7LPPdPkK7YxeGxD5i98sOySlPalAB1fWkdtaTJnilxaDypSW
6Ly4IZOZHOHEJOOWa4vqr/RRFrzS4/lqZkNk37GKUMzGFoki8+d9AJaIfctlqJGE
1ZV7vmfuchMXCyaCj4Ywfqp1zmfBV3+7Byo8HQeffxXCgV2MOqIndisIPbBpN8K/
WQZOZ2ACBKauAkBC608RAc4WBhwq8eKfJ9liQ0yeHyzrLRjRvuAfvh262WdnWwoL
Gbs5rYgD37vg2p27ZReBM2vo6TYwcSM7T/1dxyo7iMZVo4hUA03UeSv3VGq+ugbU
00iZgltkjR4GCQd9k96uYSHUnpMh033LCLyH0l50WkuklqwzO3z02EeB1vtcUUuf
YE+Xhiu+MMXbe2vv23Zn8LI9jbgATnkvjTJbA1qat4iP2MiRJzVG3cT4czSubJwU
7otGlrjuJiE7X/f1pFnAUeMm6tUBdMn0QOwSAOX/WPLiXsLGACid3s0e1O8V8JiQ
aYuIa3NhfWy1UgPw7H7K+U1LaRqByZrcIfaUPA2Ldgt86iknqyEoKW1d0eGNEKyA
XKMFN7yTjqYjMZKnx3DU3sZ8lp6YD4JgqXAW3l456XTa11kS8dhjhjE7RGGhtLbr
CJl0J/v/ihBGhFf23goy20QaCtFQfjGBoMVhIWGJuHYdoJNUMW10NtTw1Uz8VcOy
KYMctozmZiGEjg5dzAGikXt3xRU8S47XpXP7/lQAuYNOvnpvhbNfo5az4kfJ61Oy
VL2rwpXI2RAmTv5dF5zY2hiP2C3N6cjOsQUOZVQSzM7bQTLLJ21b/3QA4KS6yfiq
IEjWe9zih8xnilTvEgYCOnFYWpBt4akZQS/myRXS6/cOunQJhBCnfmYOj6s2l9sO
PshYVtgSWL1UpiXhjQ1lsEV395LLY5SxHHBv+avDhXLvF5IobDnFFkW/hS4p6XvG
pC3+5/tVkubDY2C1JxihcL5WFul5jfky3AiM64+v16DayzlAED6xpDNCkeXuh9fJ
iZs6BUXmkZm7hFoqWnlaYNDBlVnvL2mhLkXq5YR7gXYbysWE8bKrznrlObVtVMsc
KepJe1ptF9ycxzZbU2fRzAeO5n0uBQQ/5KMY2lYK8MFIuS/xTdnZiCoYU2kye+me
5+RbeKZYzTOZSfZZAAxOQo3WXVSYzjMmgpX3bF/xW6Lrj8bB3fwoPbIGvyox+xYH
MyePU2/MjI4VFcrPBYPGMNWvNVxNpGsyhYHbnwri5oElcYaZGex1kPckMc4HSI3v
jX+zbgPN3DEwOBE8XrSTaZK/OYBav+4ZouoAwcJmD9JPT6K05kt5EbaWezQoNUGr
uch1uJpPiu42cXhwL0il4zzeyvHWDU3akBU1Oi4LYW2pCkc2AxfphWGd/LYsylsI
s7Bz3Y4fo5VeVJMI130K1isr6mTdLpFnu5sk1mZjE0G85KDuYEbXe05NocKSb6sj
TGyLGZlFn1Cn5TC9CNsAQb5SFY/I4SUU4Qw6CGueJ/RyLf9XL6A6hTo6OmtlRU1U
kZELVwTDyefXbQBFgIAFtXFuP6WUU+Dhm1cDZRku35dFduscH2RDltZYKar8LM4A
SXB/4gHvSAAqS+RmWj7DeTbk1LsQjN612W7goLJZwv7CJY3Nq1/6d+gV8NVCbVib
rsy3X54LOPvDO0UphniOiHovQoDHJJcdCmv3eS68WfzA94fUJMYCCehxV1J1ehAX
g8tWvvecfZFr29VWNLvoYjn93+wwt7y/Y+S0lBGxOR+ecIuf9Nd/8XKJV1LG5VQ7
izBF6G5J2PFBeNTPGGZuOZDac9fyr6ZPi4YqtNHSydmaDUCl5ouwYSnEwnUkXd5+
ZGWaovdMdNxasr30m+o1+pWv28lrQCnkuVvXtqO2OXJx1RJwDOf/2pdUR5EKX5Dv
QAN3s3aykrt5wxpvzx9z2+15Ci53K9vElhHstntD0p8sDixPQQPlOnOtuaurzat9
6DLSlzQGIrQ0CAQp6u8HjFHycmQfY+aYcU/kMiEsgOBHAD9wG7v8hP/fjmQUioyX
sOkxwJfaBo5kW3ukg48aqxNoO/yRLev2u1D1oqzeudACyEIAU5PdyWG16/+SXTit
/MUBlw2o4jxgwl1xMoKZLORSx2beHnOpNN5obaa77F6w7/DJdviEXw2q/QVboXAO
SPWMvdsORo7Be3rPpU9Ixjn8wcZnO/7AEnpHBmcY9TOP5HAJq2glBf2BJalcVxQT
3ulKbMRAimEly+4Ewvuk6IRJmGey1Nho5O8V3SL7PmnkH56HepyL/eVBkKuphmbm
752OYNT+F+CvJCq/A5GfNtn4J4y+q0+qurjBCARJEAqtokpQxz63FV62wsg+nVW8
PoKUr8LdlKfAhQk1vyOyyO0k62lTow0OFPxgDuscwwApFf3Fu6zQ91GA6PHnzGYE
OR0m5HQocmDMJrVrnZYoQpOiA+qP4apsYux9GF7R+joHlmhyZyyAFQlB60gS52A2
OzCHPoEw5sYjQnFAqSCHhib+2NbxylRmEbC7ysXYAc7BqKwlksu5TuGxq75WGuY0
T0WSo0AenhikXamZM0XpMNUe0/tM2ziacZF3d4xpP+3bC/IhWXxgFrDIL3qFBLrJ
LkYShfTIgszxYt2ldlWsW3ajM+lkxb0IennToEoufdaV1bXN3CBqRJwqPtJ+exYC
yWaa1EkjqBV8vt0Ra9wvHx3+uRtrknIcG2lawP1aMwobu7pkp+a6b0WTPwBOL5Z8
qX8lQD71vnXvFRs6Gvg+wTm4Bnglt0GKXOok2dkp+iaEx44sTRLGlrjG91RGX2nL
xlSU+7/dYUCMowKTbpf3ql0NwCYfVpBDLCJFzCKZWJ4mSbzUK/dkxTDHz+igGtA/
JpXHSxSsdrLW2m3L9aXFxbIW9loZr2QAPsOzsqbABoMDEdRd2cGw7nmkVNy3EhnA
8LU3XlMp0+/8u7FCjm4Wp3hWl7jrMx6Nr61mGI6+8xLgiviUba3SZJKw4hFLzZY3
Xosfg9BipMP40Sg994H/tVkA0SmjjsOphtEZJw2yI/LNVkjnJsLd6HRMWxT3r4lo
jQj3tdOk1C8FRQDJl/NKt2EJBZ3Am9WlUsjw/nXvMddFPw4MYuRqhmXRDtVPc8lG
M87kBag+MF5jKLp4q64u2QqmADOB81lwog+J5XoRZGrt8Oh2DDKZrXgGz6L77SHk
8oZk3uka+nOg8S2XafFiI4E+koF4V9qShFYnJp9Usz1XsStjUK+pML5T9SmiP1zR
KM9PbeY5n9LI9EA679gd9PCe5pe7oolHl0CxkCXNchDD0Ua71coKWr8RdQUWmsg9
urvacAXBs6MWUGzKiwzy22Bri3Mbq944mRC+5Etn4+Rg9he5SW/Qrx+KdBrU601Y
fQIbT65OYZJfuoG4vtis1T1O3cjgSH5+5pjPxw8EMzttA9AyoJZtBEn0+c7aG8Ks
OXh+TIu4fwFAei72tI6ZkS8V3FKDD9du2qoFpFihXK0Ek3MTMDB5NPVvTAsEUI72
y8sdLg/+U8+sxFXkRGyL3F2luIIxecFU4d2Oxsd0wxuXeCXpuZEbG+Rd39JiVaSC
Pt812cMJNhoZk3yoZbDlKWMVmigz4rHuOhFrBm+rJdhKfaNFccsnBYX3Thxa85X7
2W+kvdMCr6nw++Ni80YPN3jg5SHw4WQarazeba+0Ic76jdp0tKSG2koCcCDlAbM3
umEeVXdwQh+ppDFoZQPqPcuZ5E8Lkzigu3ma+ztC+TN+59hPyAKDA/nx4YgAJQr8
l9qvJrFGjdpI/Khj+ybLICiPGDz1KT3aT7jeUsRxabeyggDcEggUjhn6Hi/nYHOa
ghz73ZrVeMlIo3nHzLP5tmBUWmKqNgRl4i7OYpv2yPJMqO5xkWI27jl7b87Znoul
wdyHPoH2RbqlXR6SPA1eA5/R8a83vHmaQdtnm4alvjWrozdEdMLWneM/j1A3aWp+
GsIhVK45xM/iJc4gqfl3gQ9zoHhSzcRmBzUIuEOwr/Mz80zdhyYtY4QlYq0e2qTn
ISgiD7iHHsQzZ0MHjqMxq6rVHxNqSHYuS5Ht3n77WFOg5BYGkm1vPEm+LI/0ENMf
8ZGPcVCj5OyGz2bGgljgF2gYca5WeA+Izpzh+I1H+kgn7Q8ruhnNHas/1DdARqpb
HuTm0ILXT7fPPuv6oQbiFfE1Ru+i6EcjPtmh84FeFf0WS2RWvg7Bx1mmSJOI3m9l
mmOrPocIGQuB1u871BqpsyogvDGdU4K+NEXY0RKW6CDNiitE+nQzobxMtcVXr+5j
1em7oHvsFAiwxOl2F4xTTEGi6Xvpz3jRyeJSND5hWCrjwd/HZQquQKPzWVQVjQpE
lau4BLtuojrTO9z8SaS/STuivdY7NlI9KSrQ9t1X9S20+sUbDb0lyahWKBwvu5Fj
2WvfqHnfHTbP8IZjwUJG1rG3sa4rDbGlNdlZxFUoxcYBAvKL65sdHvasT/uv+8Oj
x4y2skp2F9OwMeGnHYHXehn1C/+Afzlqxjbm+ddFA+htSyEvudqgyyni8DvcjK27
+wqLscCT/qIIt2wwlgjUQfXUi8+m85PrYJvFBkt9Yjle5wegcWWXUnNcnRjI2Rc5
cumGTbvIMkTtdMmi+oH+z2DMYTjZEvWXFytX7b2d7Ye3xnD77bRBO6PG4cK0hLUU
G6il1rxbRniXpNmnEBadqk41xSpJqdzuATVx7+BXOoyMe46rORun1LMOtcwLpqTc
pN5KI3lHsWPkBlwLkGMGKuInSB46YwtelTYUkDOUZsbQZ0QqyZ8DMbF5y9gkj6sg
E81C1nnoHZG+SAllDrep23Kc7mRpYdgo5UOD84D5+QTWqFgUSltVnRKh95qEzvQ/
NKasff8yUWriUVVCoykiZ+bTKveVp53ESMUy5i1YX1HvgSF80N4ICSJ7d4vYK5Jh
DUU4pEQjHXggDdytYuJJc8ged69fXGdRtxjFTITySieza/DPjyFJQEhra6CiwmLq
/ua6DqQdaJTm/guZjdxbgzkBS6jdL9nvdXnGLv2HU/AuYaqJTQugKTX4QG0fd1E1
vHvWer5SCM5w5PL2pmOu+NIp5gG8oXaJpXMAm9OmJDof6dSpKIWyivAoLVXS6jD7
VbKfSYl7XzF76D7LU7zPWylSLekLyhc7osOWmSM+BcOxcaqHbtY1RVERzJNQUnpF
O2RXKZeTzIMLSen2oIcFOht+TgvES0PLe+zWS7pPrsmai5DSIDxFVg+AL/3MR4Rh
Wy1Yn9ksg+8CKfff5bX01L4KGeFmDClyltO1MzVaJ23k3WCpRL8dj1PdH3beI8Jw
VzvpWjrXNF/idYC5K40huCRXJOaWTKK52C4J9M9QY6q5a18lId5QXqamBPvZZklS
d5XrAa/GHFEwgV7qMNCYz36bL53CLYVcjFRS+XDjUunIC7FsWzPralBQhbd1YlF3
45SZvgiJDBZeaI3X3f+KruBxfp2+VEc+s++SdH3gNgb6+S4nutvjEHPySyo4Uvr4
TxzcvfnUhVK6gNbME0+KAHEv75rfyqnjAU0554iRbJzVWcZxttU54Dyx3Ky5uAIK
zqsGPqfYUmtpsVAhy2SHzaAgn1ww/k2BN/UwsgQ+xrVRxeeuQm7DPCfTvhN/Vbi2
/V/6SdCBFI6eTqdoA0IirnoD/+izp9lNGnd75do2TSNmUgyiVtNXKqZs4nZV2IVt
wllgMJp8dKEj9Qqik3BVDtMYYFFf0BKQJPIze3A89+LdGsH7uoKuQeM1U6XlcTCR
3nMSULHyY+YbWXXjXSFpacDBr5LG70VgZT/Bir+3hkvT9ObpWQJOOnMvFF1npkeU
x14nes33eU13+jHFrjfP3/4s5GLeBs5sqnbvdGKOHhZHlwEreNi3oQ762mPIvO5G
8Z1PraxSlvSfacb7RQhqbf97/eVaicfXQn2M0dF2efKExPRByCmnV02897SMBVEK
POwC5O+1vJDQNKq1ONPvqL8xVoJQgT7t69W/ue0SqcT2q2n0H4tFL+5hUh9ZEM3m
3nhM5GkerKWZkFjN7Gt/L7P8+7qvr1YI+OBZDXxPsbZcI3LIzdWXxhSI53VpT5Us
3Z+0SeFVXqAegC8NRt+S9qiPUL7bpwXc8GD5TZpccBMLnxCT3CbXXWc/f1sRlO7e
ItlrrSkQzRGnSyUmYQyMDBRyLyNl9NuFXVvuzjqdhdrl8F1WlrRKW6Wo26FxaNr0
0qCle+aNjE5zn25vvWLoK4HW9njF30s96CR9OznD2eakC6lCNap7btmjdJLZsLIh
WoCKE5yODvwOvk4pyOHaS5caGmI8qbBGMOht1FGsYqfcIsotRMi/bCj67P5pUYMN
g/mhMCde3ub5sNMvAlgTrYwOwB5dRAOC+z6lhdDeDINdevR5HsAL2n9llQX66b5F
vBc+3ePu9d1Ezt+fcHw61/C53mVQ7n18IS2bARdQiSXITT4I6A8/QrR8ZjdqzBur
lHIqxa7RIjejWFzQwiXeS6nreP0gRTuH6vkKZzgwKHXIv0Ny0oYiQEl1v0+Afiwc
7FAM19FEebNUHwD+aILzy2OMza6RyD+ApvGk7zWTOEgEEZDcEChnQx4SjTIlWzKZ
bbLSSXNn8uGalo7qLg5OQ0oU4Rq3P7Y+qHvjIuTTTtIfS4JMExwYLuRa8p32ryis
AzdrEFa7Ow8GwXBEbtmLFK3SKsQC9Sstdp/NtTR3uVf6a2HwzRu8sOab4/4MJzjw
LGshXvQ9f700x44m/7ylwbRpuZpqvPcwaSCoqjc0YJIMLZPbZdnIcAgUqi7IKlEa
l0t1N5cSCaCRpwrFdq/SmhpcKIJWz2oKfZkbpXIRxZW5F7thDu+Q9ESlUIDvWQXK
WvWWko3oNnQl16egm/YnGT1e0x+gGFOEy5AqXB1AFRKPl+lbMY3KBPPyuYCAqRWS
JShknYUfPaL1wWzGlHrEyWuExdzVZKqNh9Sj8qg4WzrACAIp0pah0+LP1XOfsdlg
m2mPanGuFD4qkbWlr9jxbN3pr6+guYp0k2SrvxcA9lqyD9sAzB4fvVlI1qXLB7MI
4eY6A1tLC0aBdy2dcZUN/1od8FFqrgZmtHSYXcQzHafpyYGk/Lgdx0UHoN5qSu8L
vH8wvaOmQgsweDpTeF20S9anJUCM4QX0EQjrc9dN13u8misqi+MMtDu+xBOtnH7B
h5Jpe359YlQMNGsXO+jzXPqd/LzquNieTlpsQZ1FHxPGeedwwhjgbEdyIDPoIZHA
p9CmBGgagkDfH795uuw+AYTQnlyqC671QAmCX+f3HyMo+KpT4DgzR44jOi+i6wte
Ihvo1mEsy3yWmSPcZ5kAE5roO+cCo6EN5sRLZ6QNE3S6BGkP0UdH9FBR9APji4pk
yX2gce8mb7tHYISLkNPXa9KzsY96ow6q/xZqFbxuHY+PgaelbaqNqzG3ezS48/IJ
MzglL29FK/jh3Yc0Ta5/B4xYHWurPC6YDwQ8/b1sqb9Valcf+YzZacQnXCRaEXpy
Y2wWQPSGY6JjNJVVOcv3+pV4ww4Dx7dQzLvlQbzDidauc0vnTNBwfZIRuH7xrMpC
Ylyn/Yj0ZoUWvhZGSH9ZNPyKAUgoLk17UytSUnrgZRk/XdqKuvCosqAcZG0BcAzG
ltgORPeENcndoYGu360WhBs6xrTkvZZlAJU6jjS5JINp+md2+i9srk3sToKfy5mM
CwP4SBQ61UkicwTrmre9yFydkfRt4KbW5isXUa0HUE4A1S3XjWQCu7RtV6ikO/90
SdqI6p74UD1OBrakucglYL1IJNDx8765h3WFkBaZVoCgN4CAKlc5QIfp6chzwGsT
g3JWjb+0OYlj8bWbdpgmfYWP6hMINkHw3KhO0rGE2DPsLtqzjtl4YWDvIuxg8QlC
u5Ty2+F2zVCEZ4JD6BDMKaU1ty/f30L129JCS+IoznqtHh2gXSJes5vziLZgNr1X
MhCwllolJG/IsNEKvtM6g0UwuCB4bb2Neq/rN4v7jA8UNBRmNf8YBT7MICc14g5n
laAmG28tHosVcRtC1SA4JijbaMQWTckH53cwdKUifptKw8Q8JaaQUUvyoZMAEAQY
98UhRmvVfrb686DLp0HILso1EaqfU5s8xAAvz+qhRx6K/BdkyHB5b56pU1T5yv24
ClwGvI6EAeeQENWH/xENUfeYX4tSiEdnjb3iGOK6nsNfavqI1MVEHiEXTMM06nhP
+p4vDlQYfprcm1MeIJRWMXgDAWKDMKpfrO24WNvqyQ6N/92VocWSnHAmhlT9t66N
eOCQyeo0DrZBMTWtfE1tNUMGLCENFVP2O8qg+/Xnt7V0FqtAno9DMrtavSC6j7mD
HwX23bKoG3paRMB45Ejz3V3FGfADaOtYAt4bd3ZYjehVkTYPCFW50FwfJnyKsbh1
VVnVf3XywRmJ6sVt2N8uRv12dho84r3Mz7VE+n5HA3+kHTFIx8nnbwUgqeDZQ/lY
OE8+5GvsS6RjDg2CO8kB83KoiO1u7lOty8xT7SFY6DM281xVw3wXpe+sx80yryC0
1TbeLX8P8A6D3ZG2KucHbVdWYjolafpUDNQ8FxSjbJ1PSbIvWP60NTk+fOZaaMfR
1buqgjpIlFIpLe2yzgyEy9dRaOlyZNZV330a2u4nnd97TCePCtuRId7OAFL0uuLH
lIyQR1q9mec8WQbMBRYkVqDGVVMh+t0QL/6V9Jn9ci65NswYJPITmxVthiBE4ekO
4HSrwHBQaNx/xuAKapaMS9QwmJ9/kImCbrnR/8ebEdi8XbS5mm/mnDNZDqZSpym/
ES7dCi1FHyjCPRg9JdxRSGGMg9rQq2BL95tlI/6VppGjUA8YRaziHfgdaqsPryKz
EF7AtiEx8ITj+MyDLKFlnuGVYtjvAIlQAKbcmXtSyzGtdIFuGnO05DDF2EF41anB
oezEh9dMgMnQmR1AmfC74sy7y7iez2wOhv4K/KCpjEqKIy+cwLIblYReo7ppukkj
+Bl7fCbGymlGgrYLGrmIdcsuajf6Nsk7ydPhnjp86FGqvtQbNcTvPJq/59+iLZv5
jSZdQcWsOFqp/qpz8gx8iZHzmRHrF9d74B7ahKIeGO0IzqOnVNJbS1DPd0Q1f/AL
0aHJkUx+CaC27btblrNn6ZGq1/6Id/i3VtdnNAjlH8KjqAa5gmXMxJd5mRQ/TWDV
ptVqrpmBMBeb1obMTDgUySKsYMUsC+Qkt938zN4wOAMEeGR1al9hMyXw3FkBesLn
21i/7zHBCsE1WzXKRAjPiYWVtxYA1WTFimYbyrUl9VCku9qC04H1W1HNeAcZdfBG
PcqL7YQSMGPPAf7K7lqq5c6J2wIR8t4Zq68ldmPEwHAPURzR/vJvvAfdJNak9C6U
+UYkeULdnfE03neOJ06cEVJ7dNmA+Afo3KrpAvhZx5SZgShY1d1g7f3JLcp/VD0l
7HEqla/YCc8Wuu2TtK3kq7R1PO778EoYn0fZFUKyfbU6aYrzGu5iwsEeNgDeJaOs
spLFMFhS941whweRyHMy99H+yurJlF7qivprkpmVspBaqimYJ65VzVNWdrOxpH/H
oDACCWIAfWg3ZTOMxbXBkQzmRjPsK2yj1qgvo1Zxmvwl7bcDx2kVvEJqKJI3L3DQ
x7tdowSXvjDzubXfuJLtYJ+psjf5RPk0WODnGcJDDPsBlpYCpOzm4dkALNzB1L9W
8RfkvFKCTdi2xIvarmAHsT40pzmMRMv+E2fYejZGmGSdO5gKyFSmH80ZrHH0QDqu
AMSGyick0GJOON5D8XnCuSRpaviIA0uScHCmPQ7DvHjq4/mWojr9U2Q/MNFJ/TUW
iO5uns+eUNVCCQalN3Qz2SDZ4+cbtvAzBP3OXK/p+6PdYTbU4E0LloUzsoZAvuVL
orwBYIsmXco+GohceIIffL3xS/odJz+j+bDD/r+p3BzYRWmCLpHtSDZyOxupplml
P0cLw3K02plh00SZhu+/Fodojgk8fRH0aoKq0zkds+zqrwT2Bk3jgu6W8Z7b17Xd
AvzbcZzpAvwVq/3qLp+qzwXEq6m1MdvsozgjHymwFPNwHjcDOTqkNO2U2GNGW2l+
zNCkP+rpqud77SvpMaC3erqaugsnfMRn7bzn1GTCEGeXpAqA6ddnJPcK10IlLuBO
NQGNNaGis+GVix1CLjPjNtiEyRpYocmwckSzBXLhWcLhKZOkpXXLRKsTm60mUMb2
NLI0fLZakjnZHQdMilwCRZihbcK4n28DyqClr6MTDDNZnLNMM/mpY445GRLyZI7H
WyO5SiwXP8EBSGvwN/rrCx0C01TLHWb7o2c47bB5P5b0nG5kI4lRGm5o7hqqdfer
bhlqQe70lvE+HNRNsgnc10+QIppBUmbgjYRLB1eCkZtSXVsM0IldZqLkSKCvdqFe
jY7H8HyD3bzU/N71d0oMOLY85chlgPViHns81hxSgxy117e4MR7uP4y4R6KTkmF1
7oYjMIOZoipR8x9GORRRD6s3vwSvhYmIbC2hrqXoJ4m6y2cSwSz2qLVQwINM9NFH
vYynDzwqQrnFqfLphtHafcGqG9Q1GAJHFcuYJFInvzU7EqOX2IHgL98Czb82z7E6
wA55Cm4jMLIKR00ZEo1cQO8iTWeyOgxJwiF+h0cYpVLqzD+JLhDjkbclT3xEoFph
3J+cNLOT295/KpsJRO/wEfeKcSXHP2RtAqwyT+YRA4UNuPfESWHUMFOxawmak16p
/rgLcXrQuMjPDlmyyFibC9Xc1TLWUwBPL8EVnAWDFskvb1k2YsruZWD8LcTKGQD4
1tqLk4euk858aoReGDZlzDNEHM4ZtwTRYU2HAYRBZLZIMlfFnjoykCt5MKfvscjr
5DimeQnWamH7ITlTgg67iRIrZlgf4zpalzBNBdcMIZrpFInXcxFPEOocB6k/SYWe
PzvWZp7vsjHMV00UorJpUjnB15ZTeABvdyhyN7nbq3q8bR3o91yqBCL+7soxXBfC
7/HZY0fsv5WY/SKzaDYDmSDgGgsjZ21hTrp6IUusrR4y8ogqJ+UTESZ5F9mr6lWY
xmpLqS2+mAslPWFu3YfCSVdiE1cyToIJjX2IeXBi3bwXWsrTzjhoWVTaLDL6LsX2
tOdekBq9vhs1H9TZ8j60gOrsk2Xti2hiR0Bry0twz0xQ+h4gKk/45A7ewpprmnYN
UF9rifbP8aCyFiXIAe4N9dctY57P7Ht9gw9HB4sFi+TVcWmUxH2ZsTeLIG4YFoQ7
z3tw4Lv33O+lqr6mlkjOo1Gz7Xix1OzdZffUQM7rAG/TMuyMFKgUZRMirPcWKMVm
2DgEes0Jr13qtkvQcdtlYfwfwcTXggeImbfGZ13y7/tm+jwhJd+NhNAsRe/tN9Jx
FxnfpyjL3ysuFWsGoTgBQp14SvpBE66Ak+0PkU6vsWmhMGLaNq6/W/rtorcF8VBD
HWgtcEdalY9aECD2HJtMoCuluFqrHCMXcPZw5AwpAXjOnYZ48syFSR6xO3vnetC4
9e3CzCi5PP53hwmigjm4PTXw6mWv4KfyWnIWYBWvom4Sqf6IQa6PYQTllE72IG1S
QOLsZUlLL6kbXTLbS0B046bU22HoIEPQcYZs83mrPzKGrPKK+w1EFGiFhqn9eESc
zmWnUXYs3KTttJAgFVFH5pSBCIIpqyVmrtlFkaJ9oxsIf30U9zSR8VMVBZVlnUrv
Bx03Mqd0R8CS1BXRmfpcMqGQzn/yBjOY8SeesSH/L3pUIhHjd57TFLb2+A7c7V0W
es3Zj1WJi8L4ARlfFMkn5YWuwNnfeHQOk75pkSOppQ0XNdtzkQ+nfMokPuv0mC3O
2Mn3LIAAJHiHmz6l4cuQsVt56HujOQEIH9zCwjNZEqX+va03OLHJMCezCeEbh6H5
e7YNNkMQGZf9a8NKP85ulcMzANjn+zmO+HIXU8Ln1bjwd0hGyJTD52m8wvYLzY0y
Ryv1aQFqSS8dc4BuXYI4OGiZfzcRTJPfJpEYy/GIqbp7w4fVOoTrHCYEseupjZhQ
O4FAkjbP6xfkRFcqmPMv42CWWClXhy2wdtN1mbySl5ulPlw/7rsVplbzjpuEQdRI
wXq0dwPmugKc93FlPslWGeXXRugZGLZjmjoYgZzmwiQM0zMdK7H1g8L+BN1N5GbL
h9FbDRM82seoIuO1ntdoTjlhVJYrmiYYbsjGYjg7PMff2OaNh/NIZJ05bA/3o44Y
S23wJOPZEU5ee+fMw2h63HaF6zTuV9O1NlaRTtB8zDcKZRUoBMsNE2Kz50engzwd
VtDqyfpFpYn7o8Fs1RJnrkVm58A0/xy+o+qE6SuUnOEB7xr06bU2PEh/KmM+NnhA
M38flpR4/Cp5GgMPFG8R/ZiSHOLbRd7H48QShObYWNM4EM4A/VcjF/5Dk2Tdu92u
OZB1f/JQtvQHWEgYGrxqS3yIdPWCv/DvVvxD0ECt2xVh8RpPO9q/JRekVzFQh2GI
xuzXjzXZGrXX1aT9PqI7Lg9mAZHFLsv90t6/7BuZYOvUKWGcdo3PdXI5FP65mXRr
JFDzGgqoBmiGUfoY1Z3krDpjqT6qTTUR/iT5wn4T+ack6z1Q0fnbZnFROPCvC2lW
Lztwq1J4iQ0d3csyI9fO4Vh4ioSlkzpOfwXghmFrwM8t/aELgrEr06IPbyAZ0/9R
RdJ9jHiwf/z0Ocxlt7LZ3+Kf7+8jZqY+zV8v9ElhaACuB2/jT2w29K8qhx5+Tcf/
Rd831XJ9HmQaW+JYGboTgOhO0sEjc6y2xDca9JPyTIWUgzyIX/MDqeAJsflhFhIm
gSGQ1p+WLaor3x4shBHrwdwtq/Pzs23cG0gXefEQmNwK65x6Rz6GgLyFk/t/kMfK
oniOZ4l/o2ke3ufuEwZNMuDTS45AgywjYo7iAoJHTAIsXx/QZ0/I2y75ca/1c5kS
Xo7noYAg8A4OXkXIreMdhBkBNRZpZgZEZDsLKGzT8fbez/tWbVU3biK8/+wUYAOy
DWm7qvuYcYGHA+H+s+Fgbp2P9vX6gheXK7sXU9uA7LYfXygEyRaBatkaaud2da/s
H29Vu/km/Hj2BbZqCtKiQes6+3Ri/Hl0ZzZUVbZcHWjvyJ59UErhXhAkvZ5NC9dD
7WCMKoj3X4Nnc1I/anDKEly1wTgp8YFcJnL7pbHG9USJjVGhhP9ZMw1WsUHinYVG
+hYl12R7xqkn1as+whsDUztoi5J4/r1JsbMoptQt7HYdnngaa3L21rDemQb0QGYq
k4JHFaz0D2K3FAb/hxODI7nCPH6CO3Ptujd9rDPSgCH5tXmNRm5hRsR8dtkRmmEM
PFNjV5FIipui2sgkVFSelnUoLNFQXrkuFCQBw3tamnrwswU7IBRuh4CI4BRZt48D
pYN7SR7gJgJWRmUAe5d1ZSHYuwR45OD+vRrrTrkur+GG5ua4sN5mroV1D2U6IanW
lc9GG2sLXOgzH4+3IcgAl/XkNHNjCxI+nQGktpuG67TUR3vZNRThEnlnzwdmtM7G
eAteIeTkzMsFqkah7i7IXzbFC2t/pW9Ul7kbZCS/ioQE4mu+Xou5hqOHGbk6Ie2/
fw9+LzUjwAR9seAXbPEmhlvxbFYJBZtt/XXZmCiLS97kx+QsL12o9gNLhyP0sIoD
erp2nACZL2avAmaYgR/WpAX/deKCQhd44Y8S0wPGZszGB+q4ir1NacdqxnhLvjpM
E0U028cUYukx1B7+a5QMKyzXtbkBBcgg9ZPukxEb7T2e3Liaz7Q0O4Lltr65yCrO
rRQMKvquNav6LGnaW/8YUMTB2f9SEArqy/tde9o2oXbzR3IZ70jfi4t6dzRJVvlA
uwxmBctKrgd5V+/u0HFkQ8zrJ3eeuX/INA7cn7kJpyRmMdq3cM85XolP2D3PiNA3
LteNPH3/0k47cl5bFufJxTKQTdvqEkc74DWxBro1fymfkw2z2Zu+QPtIluKov0Iz
zYb1LVHmuYVNaNS2B7tEWIxpxa1xVVSSiUwPnYtLQp4X8HhJ5jl96iYQW8aG1/BW
PW7zDtYYd5ZSPHWXCbrUAOXdiwGRHvljiFCOE1AHhe1Hkg6RtRYKEZgM371wCoab
gsM6LJo6EHT/7Y9tvurPBadob/NGH3wufVFGs94SlauExReraF5F++yO5BpUsBh+
SRi7QkfMdsuhN63DJ3RxVhUFgsfgKdvqJNJLvfDiLpfKgYZSEMqU54OCDu2e36zt
Btfo/Br7H5k2P5Xo2DD/K5G7sOtDVWnKT9hR31x5LBghF624Q+1A/axaBpJPBY8b
adML826zbPuqxA848wpfjgFL/RKH6WoeI7oKVePkY14A2ODNpyjX/83lxNr6K/Fx
ZZ0iyIm5X9VneKPK0b/ILHvJp7a7krTf810D5ajbc0AkR+zagyd2wCXBwr8eforC
vy4S6uggdK23ybbljrPTYQU8831SMNtEIHVYEldaCY9sBNl8dvWGR9+q1trNMWhG
TxMpR+xFmAflK6eB2XtUS0stOuF2Y1REtBsEK5jypgF7bIlEcooG2v7et+2hyWKS
wjUgb1sinowJdl/UZS+QZ+WlnM2dtQVp5G/J/3xjQkxJS7UMgBl4Rh9zS4ibBiLo
4dIp+CuAx69HHAUOsdM3o9ncsstkEceV/6QLMFEYZH7hYTe6TG8ifge7b1vJ6fq+
BuWcOA3QSdbEyX4d/HnLPOZ/4O9GoVah+HxQDveY58UnqR4QLC3N/6zeG06z1iBC
fY6RTkyDfr/5WkX+f6GvGbgcGq5g4O775V1MkQygZDyc1jrknahN64dkXM2kQpSH
KAAuX+w3IqXpB6HbNedrHEHDb+vdUkn+JvE5eooqzXzNUVqHlTsutj2G0767IzBL
CcPv4afM2k27NdiGPmkIaHC0bHteIfCuTzh0PHE2IItw7ioJGYMfREuWrGC7GC70
Lz2BP3KXALSb9JtiMdEcvbATCW2Yenv7HRWj9c8zdyXplbUoOyuONnNIfaqpIPgU
RiQ6fwiKpt6AgJyWHYHl63Cb6SPuDqjt/fwIAU9h5Lh9x09r54A1FRwFdYoFTG4j
c1e8oCCH/x9SmlM3nLMziGRRf3YPqR9qcLGUvZ/JQyMnIK1FwZe8r9PPGcmtdUGC
08gtBKYEA8von8fIEewpOj4M7LYnBPLcjMNE13sPLkqbPBiI793tNMxrHUP0Z3v8
JAhHvLCJim5sT5j7uRV63PLB7sYxGKfrW1dXAQWXdkKkr3V8CCxkithLPksIr2V8
tJGs7yWmMdMz3qzkXsUMsnIdC+z4NDj7zNVKMig36h6u6n+opVscdrjdkAoG2ONA
+uOnVIcuY87yvpEvo/fDV/oO1Wt/LJKyb5XWXjVO/j/YIK5dauRu7jXBdgvJjMmC
lN/biLBOq8d2N0RriZW8gjhkFaddgdgBLwcyZ17whuObFB3TLDJw7X20G8/J8mDz
0eTzMihTcFxd+IYONkgy5Dj4GBGeSMU8mkuVlbV+evvz68Kywniunoi8YBtswB2O
I8aDnsgbYnjVgMa866T4Ajbwdkn+cJDn6prSxpzGQ7kpOUJaIYP/hvm23LEfTD/e
fMIYMG0So0JR4Ndx4c8x/PNB0R5k4SlZxegURTsT+Q9DjrG5hz2culI0tGf4tnid
9vnOydcXTAGcNhYNffyNwplWEiqiu1q6+YBgvp6wUHbdT13zrj2zKzHv3Jssvr9u
HKdJGOmEdBQ7h96290pCQ5O47EJBnQ/sx+1mBkMCxLYmPj9SO20jAgHBlXthW/ae
RFgxFG1785VE7wcmc7YfwVjeK5wrW7mBWnRORx7ZxE1uWgDpPK6sInUIz8mTffun
/meGDTmCVY0mrtAQx0XxHBze1AA/nSsXrsWCqMtSZLKoUyDMAc82McoYincQt8jF
KfUQkgww8Geqw5hn1fdoHiTH4MuvhIlWLm/v48hE7qFsYjrfkD5oBLo9bDLRmWWc
td3OwxE2eBbz27cgsq5j/1SuaNb7xA/DS613QrvbGMx9lO3xGLmFRQYUjleV6BYv
g0OVO0mJSEYcT/i9mxG1rsmdnMgt8qRIXlUm1TuEaxlRELkJZaZz7bXIg5ke9922
tinFWf95t1Ij1N5tmKCYborj/KmSomat1xoY8N0NiLuf5JrWwLLpuaUJ7PxC9vJp
J+p42lnhGfrz+TIftNwf4r5i0Lg6OrOGQDZxfOZ/+GimQY4qY87M42cJxdcqmg0L
matNlf0FHcpQ9d0GUZs8grHJwSqf5Ol/JeOjwDi+vIAMSBICLVhEJhVSbBquBvfv
Xvjt2MdWBczyNnJXdZA9KdEoD8Iza171yek0OKtGXRC/Vhk0Nmte43knXQ7lTxi6
9ytn9Xp6iI1iI+albA2Lmrh8UC7jbgIAyWpWfnoktzShCxIdPIthMWvHu609vcbA
AduNqvlOfLkNNe1S8TY+bapx7Op7XhS7/IMj69VlyMwCZWH6AMLtYXrXPgqLVmHc
Gi0xTcx356UbK34aETqLv2nkzXXjLuKZ9Yb+hCnrIE39LWglo/VZTj9LY164JAof
JHWCbMC1/KpW5CIhz6KMIoes/ESQ21mju3Di61Q+5olbDeOgL/aoGw1UgTQT/qvm
nTLyQ7lj65w1eDOT0NSv0yUI2j3vlXNnqDC//aUAurgSp2Q7qRawKU/P2YiVKGwV
zP7HJCLdGFZGh9ayG9FnbcRNGqJeMBLJ3F0bIe6pEVSaA5ms5BMEdWCaqfMNaZ+C
DEOWSo/0fuKwDZq4SdqOMkJBO3cn4HfjSmkmyvO1ETdSLBQ/JNpbWmIe2YcjavvZ
A/RFeU84LQE7/UgF7d/sY0I7LP04ZSiAFHQu7P5EWqGIy6wR1gnV/Avxk+NK/9g9
fYZhvIDTE7Cplt1k3w1BgauNi4t20Ubrl86WThs/m/Aj6BmQpKZZO2uiMnKnaTmv
F0yIQQ4SbH4Ejkumwjeg7ti2+UOFoRb/gMyKVVwJVG+dENS5yctS0pD8z1ChoHTy
aoVGN7SnvgwjDZBRawx+WrNOQKsKk/VpiFaMMxOo+jZZ0G/DX5pHm7muqyEXFd5I
8a3u5U2J9Api5uauuoNx1PFE54FivkKwF3hFy+WHepgYU4sx7Id1pggvTW2kJ5FG
RQDR1+pjebgYb6rn6pt+tgVxqIUJGl6HrGHpn+cDC/GuPIftdbNhRL/JNw6ovbm8
BfHBGd0YGKXfI7XrL2byrRK4SwXixivabt5c0kmZZFJFq/o21R9m7B3kgD5Nvk1v
sF6qc5rVdpQS2a+VtCAUq+WX60epq0NPtWjCoq5fubrKC7b8JyJYxPJ3BADVDqbl
DboDH1Ka1oRPX8qgYGmfNnB7LugbKVSV6NKKT/z9RyDoS7nlugI2YWm42HbwUUXG
oHCSZRzB9twJIF9BmWjjaQCRp/at/tl4RT0wxk5cWOGyPEY7diSOUnRLV3Cb+zDr
qIv4Vqe8zjKLvbw8SBbSePSG9kl1T0nvqXd8D36an3ZqVn4fplWPJDm4ye4IO+WN
hTjHQnQZStzJFWcdeijuT+0iRIW9Z5lkr/d4qW+TGONwfT6s75nXYzyjBBtt532B
nfd0ku8wtaPpJd6JoE1jK16t7dSoxmrKzz1SQp7WBwlMhq0WtUIL04ejwo9aKodn
/9DKXzGoSmE/CK9T1Co0+C32e/smhfi7GSM6Szvr1Es1WIgLFrcKtRDcReuRHIKB
wOKoBR1sRsCKZX4VilSpiSDpd69YE02aO1DijD5o1D90fXPRFZT0A7ciuus4oFzj
iqAZ8I7HBTJetWgT8MyCCJHdWEUQ3u/3c8gLKD6ChaKW+sp9twqquvxbZd09ud6C
qbuOU/2ecP4TIsteetyrlM1cMYapo7mM1JJPpOvKNl7UEkIV6xFW1DoamnMp/+Sq
CLtekT8ydgTcsxdhznU+DpGqK6GRHWPUFmmHLpYrT4swylWRe+zfkEoVGmzqbmuD
j+QVuors9CLYILPAMYhK7ZeYTKnR9/zuBXQIUNslKORL4b+iAijNfdCboNQzDoVi
YGAENriELsYv/cGBfsC0sUrJz6Lb9q0k2S1vzJRrU2pv0bZhMgInPPqIYrwRcg/6
U7pef+ud+KBT5b6Ri/8XlguICwdId/SFwMxo+Y/AwE9IpADQLVvaDEJSRa9IBPDd
UZFJRgA/oYljxHa+fbgzxyuFqvaWF5uQhrEO1QCPSqlNPVK7Mr96UMCBav9qR3M7
bHdipNa3JwS6Z9ZK/uUCHUQqtJrTwewFPQbhh+C9N9irICrfBrSWYJ0X6VsZtiJy
U5flp+CCp1CjWTYmdA4Uuo83gxZS2NfemyqidfcdpI7yFDBFGZLqJltIVHha/Cdk
kpAZr8LprkaNmd8ESSEqXrkJSgAiYbK7JW9NJAEHGovRy39DjBhuIO/whR+jTJmS
W8lu2BOu8hMyehlZIgr0W5bG/2NfxxhSuLYhdoRcBCbnQKNQ7PEPxpoogNhya2nj
sJpaCl7adc/ZLxds1Eb5GVCkZOVO2fQalefE2CuuLMtaLSYS/gBusd61tEaTp+Uh
IXedgd1f5Eu7fAo7fx62xdGrTdbTXcvrmnnrqIJ6J6F7BfQbMKRPyAbKfDg9uBa0
8BKXGUYXz+AqzAgMqay4nOtoqjkr1eYj7zl3cvH5TzXoa852UWpzhSsCE/H7KOGi
MXpw9PS5i7GcGZsIaaCVZWLVU4gTdVDa4dJZ9jzw9oIcUpXZp2xSi14m1X5+Pl5N
EQDPZvugdEt10GLVH3/YtViCezbLgDGaz7taVp+V5U6HwXLLvy6aJOBsA1g3M405
96FxRTydy+ZdaXa9x1uYT8EVEzFzkQKWZFRy0hyNhOP2ZApL6++9rBumulUz/LY4
ZizHAxYXq7fBNMm4yttAf3qYnLc83r7BTVM6UDIp2q8rLvBdk/obiQE/t8TPFn6E
Et4AfoW4vXQqRheslWlI6Ia96myVs8tJxxgSB0sOu5yBjvsUEkcjifp+c0NgFsDR
toEZ1kY4ejxxNQB6Yqopznjt1grKj5dRfvu84tWFIkciA1p5RPUnhJqBS7UC+B57
4WwK6YWmVvz7PmXqnyjOHRLrJQEazjWEkl49mtBGzWmol7lPnqWf3LbS0l/3IX+t
VqYyVNcob097P60wJ6u3H/H1brAOiwrzxvENccQ6JDpQTlNjzQOD5BruVClo7o+4
ykX3fygXV7EfkfgQ1mmpmgNrdi+N7s9ayWk/C556MrkEpyHW6EA9pnsN3wZfZVue
V4xqrieISgSisP9U9p4bdv+0I5Elozhqa1qjc1E3mna3tjTWAEmhyrUqsGumKc8a
JMFo43Rj8VnEm6VGke5Xh025vvZaE6s67W1vbpEFXRY/jbS95geNycqbH9hm5apt
0DoKzw3f/gvTYn7I5JFW0nb9KBRFD8H/rH7o62NI+VBk4S7PlxHJvUl5Q2yjx4TW
US2lowH9ODskhYKrfWZ9lklhj+s64A3/B1w5bQgwRRUtmJrluDeaADmd2At1J1U5
kJlCErFhG/+J+8D3dENbNMC3dQ/liLkXVMLx4X51EKc8A1jKCOwIDUp6y4gEavrc
1gtUlmhG/OhhvincV2iyKcHwmnxEUvuTZag2TCHsF13EhSLMErO1M9CWUt45L4Cn
fRk+dhsEkM4bFzWzJUY0bFJr1MB9SznbrJRItuAS8lPZ3m2khFdpzIDlP0BaD7PW
Hp+niZSaoalS+y1drimSAehgF/lHom2a++0gVRHBXDXNMueaoyGc/ObSukplVViy
EQXxI7A9ZUiFqC85PWaF30DkUZtzwGb/sisuGohaPvcThnriaiKqcRx7Heal3KJh
NVBQpDKXfU7BTZ1TKv8d4Riu5YcMaDsf+i9v/IAS6iY8Es8WYymfnYJjDNdmG4e4
ND03+u/06ugMUXndVdaYygxvxo0XWbMPHRMJ+9a+xXMivtAmAvTP/80UO7Q35aA2
nd0O48/ooKQ67ZQFiTKfJsn4dcJLWTQYYlgFGZxWXzAnpT4PMH6H0g4K9z9FgB+i
paBMoiYgnRqGLzc0iSsK01ahg9qErm6ZNlfKU5vRJLwTwlunttXUtNUL6rCEGugP
4SwrXHuliw/vyuq1/1EbERY4+SSOOFU4o98jnBZerj0BUqHBoiVQLh9Q2hFSaqXS
KYPIwXmiLSAime+4AHfFKjqRxVoAvWIdofD5WB0Yo2NV7HYGK1UM18ODoA70XHJL
HkIeXnPCsm+VBcWgCuW39nWkVfvZ/eNoiQvaJDu+fMfgqSTHi6tt0BK1wy5yHns+
zfrwxVwmkv23Gh/QCnsfYxu5H2MQlGpThtZYq+TUNthXeSjQvQKZh8/oYJE8DCAA
GczCraGxY5mMNGs+3zyLYj38x4cOobApT0sKaGu4XPyaRDWPxl2eh4EH7NO5S+vR
F+p6oBK3rqhJQVymi8Lw9SmP8qggFwnz56L3+GJm4+fOv5FUka+dgVN2UPDgnjUO
IGaXWiKHv1RfrBuygq0ojt2R9NiPGmIFACvdwQtEq+iTUdr4GhpYFg1LRtIHqm9f
pcqRl9Ki25nQ81Pc03GiEaNWkOMI927iD57bV5Wli7HmBBUnmnr4dRJQEybkLBbj
CQuhsdBdytlFDNGJG1SQ7FD+nRKuOVdv0+9JqkB4cy5jqAiGfIGTZAkOQ81YTDh4
+fuiyUUb6Gotx0UjvxhQOJNvWUZj6KxSHQ5PKXd10rBMNPyKjkJjHhv01TYEMsxY
KJGSozzOxz6K434iHO9c8XFI0j/hrJhJnnXwq3QXarlVWrRxaLo5UXP+9qcoSMN0
SBpc5JaawARoSCE8aJscvk2IdscQ0YBDD5ebs5Pw8rsDUP88pr0xBc5EZ9iylkvE
fU8Z+wTtLf3cO57046NfHF84/FYx0NiqIDZjIWgZvC/fOvA8mWGUpcN9g3DOxO8Z
G3zKnZEXQCdMALq/Jci56Mu2+oV/cvCs1G+ndLC8/5z7NZlRKBuv8VxHi3gWcG47
OmsXo66XtJEYz4964O9p2KRsuceo4SRq0AIN2N4m48vUcnpR/8sF0kJ1uS3c9Rkz
uhXPg1KhCCWTtAJrWNn5gVS+Kvz1kACv5uLKaNegApJUte3X83SpFrPHOO2SR0nJ
HikWfdtxyzg50Q2VMahOQ6qWd7+ni4MbwvqcXJEUMY4ZUDAvMnNztfnKFi/5x6y/
AusvsATt16JKfXLhk2m7UIB8crfnNqhlUcGls4G74546oM7jnDLkYL0k3JE2pfyn
C53i6frLInmQw9jSkKmtySTnc0wcu7LFM2UH0kNMCgKdtu44ns8cD9YoQq6Xyo/J
Lx9l0+FnnSbc/e7kmc6saijn6R58AR43/qIyb+xdCD1epTX3ZcGyCjmA12LCcAEp
eLYU+e1SxV0MTNo6/B9WAO3suQ3u4fPQpzaQ0Yvv3ZFvu1fClTDmUFCzJjV0PEmm
s6N94GmjnZHhRh6frOvydWTACwfQ65xBBSBd6tE8s5cZcOnZjW+XAVsJuMY6Rc91
/W1VesWy1AuDDtEP1w00yejRacJoTPqcc2SCwjCppQayf8kssgsbtC4Q+vBvLkq3
wDsAJI2D2/fJVEw7z0aIP2rFES0zSamnn4h5lCnVKro9pTBxxADgN+ejc7UIoU3g
kA3/2zcODOuzq98BlI7YavSF8jRZWw10hnTuE491Z+a7avFbUmDiqCjwfK6GeCJr
tR/i9XS9jO2W9B/vP8k2QZy5dULMHo5jpxPcKDOsWMz5bUE7I9qYODEBOwDefbrO
MUIUEzK+UpOk2+zBtw+Z6epJmKEHWsmggtOf6ZfNNGXl64k8lMBCTY1rqNE5/Cny
DNbuxJw5z5wsTVf5lWR8lQI2RdJAt+mI6c92BRicAP7NnO0G9rT6RIbFGtKq1fm6
s1pp7YsWCe3FHKHjh/x96nECFirYU2lhA0bsRgbnkqoBaLRgAxgZQJVIquGgQh+T
mXR7xxVeOzEdk2IqSQs7u677yW4X9JqoBDeQzjuNNNnKYq6sGaWyYCIF8mH+ts0l
bxTPdhMmOHK9BKzQOYO8x/o13wfTQhSmrl2UAzCB1DUf3WK40eq84BKBeZBd2G28
HMORHLM5HoFR3ua0XiSPZJn44PtHy97K6pH1vreq1LvDBRllZIsTjC2LyQPvpOMT
9Jk8de/1v43T4b7+gqQGvfs+x01HoeYu3CWd1jroHE6rP+PfqzCo/nB0ujKLUec+
sO4Y0W7AMlUXiFiZ268YziV4xU78vbEVRsBYhIaylQdfpwnm8K3fHQBitZq/OWfV
RGrzynA9kL3vLlvEpT/lunhiD6b7ig7fKWVuwspDLT1R2ZC9KCUTVUbRpyY6Utlu
9J1PjAuaaPPJ36qHj272a/zKWh8YQUR84m92Y6wiHAc5uwXJ876RUE7gI0TMQ6S8
SN35aiHgA7Lqa4S3Vo6KuJ2fMlWHfHrIpPjZUkxF3XAbkqoNR1PchDtVI/oIGIlC
sy+gLuPeOLais7njO+kzWvNqw6sHO+a6bkyRjvlexfBq5PcpJVdarBx0OmROnbak
HZlqF4oAqyHF+9hu1W0XawEd+/8kZFc5KfTZ1etH1QlRYRmzBrbOLpw1r3bRt01s
a0LPJAvhLypnlFWa1Q+xmEL7x9N/Z10WUy0xQk94xyy69fpx2hatnwz1VPidGYDa
p4qKSYZgyCFOvpFVMZppnCQwPdcoM1TU+AZoktNHJ2qED52zdnJBFZtAiTh9qh3n
Eb3CuX73woRYa6cuqpcYWAPQlYAXo9Z2utxZkBRq0YBzRp9zJjdsVvZtt+qaso1H
KneQbvi/Xe7oCyoLR5RpTkeE3Qh/yrMgagWqrXYK+vbjQo2w4KWrRCmo1a8uAWCb
62Z7febUvjOIj6v9MzEfLmgVCt77cczKBdQDLJT2CMADu6Y56UjJgA/hFRHe6q+N
F7RTblJdVM1HWhmIWgR5A7J+UWrX/K100FvYLc6aNLm0hMV9WP0DcMReK36EtRJH
AYaVVD5V6mAuddl4u8EX42IM9xiKkk0EiN+HJ2y9u9uTBKeT68e6PMwuTKEi1gRH
zkO2AcdR+fa8MlnLIYgieUsmPMEGY9hOE/+2UENq60nMiWI23rabM/8qNZBaqaPx
mv9ciXvEnlMAMtpLtO+TbmLqxuQG2bjylc7DU5n4y1BzkogptvDoFr/f+dMw2fOL
FplgyV3NjEaOpIIMyzjtGHD4dchRY/u55CrVlxdxAXChbCbn50qu8DAqje7fidlV
eK03iiUUIt9uHk/cBfss++EQjQhfoULbPdXJpTwhz4Rvo8lUB1lRSkdnzSyrImBl
bccz3DxWfy9TW7Cxqfbj1Xgw+Pa+K0ipI3Px4SjvvRViVWVv5G4dCDrYuUoiHEMt
qbCiL7wuxOgS5tyIwnpQJk/3TbHnV8d/Y9S5WoXGEDqaZdroaiu7Wn4G8HIxZTQm
2/J3jwP+nd9xhsCk1bmivtnx4c7hkvWUhb0ODzpwfObeY7nLRGRR1qkAv1qz571x
HGvH49LEc7gJSiBerZqoeYoBgj3H5UNdAowy/dDoMisI28AU8+AKLpmahKeCI+y8
JmQBWI3WHQ5I5C5ofAjUL1xxroPtZMBEPG4ljfm7XRutn3Xhkm3Tf7Dw93ktfp+w
8yYrGo/QlZTfW9PXkTmaKsG6HAvQSvj+wkNHRKWzNyAEqv1d1ve6uufHcbjR3ew0
Mtbktj/XOxrjRS0ETIFSNNoK15jdZ9xc9i20Cshkh1kyHJH387vU7r53zNxGRpLp
s/Tj8iuv6Xt7lLkBxDR9CzbaSMCGAVs90lFMsHTk6nf/sp866VYj6T71CxnYftY5
jMDlYgHkLgpT/ZQ9ZWXduYJs4CxM4ocenUtvPku5jKVOplk2ElNxW+sFUfNrV/ZI
4fzttQGhBWhcfESsaEtvqccPuUqJ/tAFfuJcMdJP7TA7C+2aOORm5/UJ6Xgc3bbs
G0nwBQYaCt2DcANrkf38nTt/Q+0WchDIgwQAJkCPp7Evqyh/YkchODwZqyvyYlZ7
c9CJyXxO+au5IbjzEziFlRvfq4tDk+9sk75d8pcZ6w335BVrfFMi52QlohjW5R21
V8GZ+1jPDzh5pkUeS35yduJZM9YzBAbiIc/3QiNIvZVUJ+nUgdJfxm6h9qufo/uP
qUuRPedBZxcu0SIUZLUBVu8haAiLKJ1RwhBfeawYqX3PC1f/r0ao215khQ2r2B2B
GZfkp+fVH/IwTk3EP5++Gww3seDXv1PHL8mRLBwavPcvHhBnIYNO6kzB1UgmI1bu
Uvgro7IqFLEx7bzBpLT1f5n9iWqyJ/pujFvRcABYr+ySVJ+iINq9Tx2jqDerLVQM
pC2iUGPnJKhbYEzRZOkyAeaBCBlYWUq28VA4qxx3TejVfMY3m0VtIVauIZoe+/fe
JiiUourVwa6qy3YhyLIB/cbl0RAKWBiW8sAbPmZzcRqr+CaUAQ+ZQS/kh09t67ta
nvfDGJXefnGFsZcKD5V1afvPw9BIDcHfcj5yyDK4Qvn/Sr2p96HQblafOt4C/PZz
qJfuvcU+aC5naq1WpZuw0ve3bVPCLGTG++Y1a1ONwf+jTsELJeRWOCxZ3PM6WOWy
IP/dTeK2C6eCvtL6QQu3PriO3RYIXYujvp0c83OgoT9djshJvNXr/VEezcH390aq
bsGTsAzINPxuDhXK1FV7/2uaoh97vBIsH1Jwycqm6ju6H3Ce6wx2TxPGM36q8xqh
fa80A2A0NYnF7/xTec08YEdB3h+wIevv9IfmXCIEnId4Ri7SalArKzl2rU01m1+t
h4YIn125pgzqk9mp2JOf+jNT+OjqDWpGaYQvOYiAoxaYqYtuSqgD+nUGC0oR7B+A
IWz3DrqPB+TnxCyVCyVrxhAbwr17vHYWFxQ9x90SLELMVU1RspLivnYGYir9Tok+
1Amo5siLrFgqALu4bXHxN2ik70cD6B/zUpdZCdFSkCGqLWf91C8QpslOXaHlp03V
iHwt8z/WiJzWMzIb+wJ18CZ00NVbuesEbozgi2Fw76MDRK9WQlL9Cc+fwMWiZMbm
VUgoRxLif1VDWUAt7X3OcS26Da3GHGbIfU/cyyuFIS3lNDPQBiU3oSsXz+s7ZJeY
rgnmiNfE1uuGDzthbPtsPgTt+FeocXlxwW7Rg1ytIRVfz2L4SkYxRivT13pvfMJ+
UQGhHDslcfxe6TXjnjYihQWVoUWJ1nwKA7kj5d9U+wBJ0OLkpsiG0nZ3/AE/mt9X
SQx4/Fr5wQxWWz7VbQf1E7GJjgpZeXOx66SnGBfpDTcFR9pWskIdG88N4S0XxoSV
k2qbNUkp4PZfI5d59Wn1KWxH56Hx1UjfJpD1bER2Ybyd4y+W2Nl4sbqrJtNjzUgz
sGQU4jxfGTV30WkWuSLOoAH3U0iS1+gpgrz53QjAjA6HzOVFEZh/xO95gvlWQCYx
rlR5PLOLibe+ZmRPiSw2FmmCAMoqy8uDMaEvhNYpCtXTH6jjhgiikoO8ZY7sh96o
qruXidMi9qZHsQkRFBrR548sj9WASHLdzgQ+/Ve0qekOUhWxd9kJUANULqkUoa6v
dhbRWr0b64Z0im9SzGpo1rnYdURwlJsbCfUnb8rO2QN9c99muMiX69h5HaBqjhH5
xRwhUjQOmNLTcG0E9/HmSFynyAJ/JEVGx9SBsXQMIYCUcgEfpoG23za1gmf/lKuf
Cvg4C9/rei1kf+l9+oDG8uScfMv2jCfzQe+VIe7K+YvzRhPl+f9WBHIuxc49Bo6F
dgGK7Ki0xwWZNr4wpFgcan1H3BY0a6O7gnWryXzl6+Dtj50PoGT5+sxJxj1ZCxbf
Ao4Bgkx8uS1Qo1qEHw+p3KFnTEDZRuYJSnDzgQEDtioSuwJxp4reO5zD9RtdA8Xr
na0h2cbXBBhJUDypn5g0+9WQLMARKo9L/PLVHnOjaIaWzC2cpQGDYCWFNh7YIH35
LwXkvtDs0zdEHFfQYuQvnCg+RI3ouYin6S1GAAPWCNaTU1fvUlvxe12sz/P7Oh7H
vmChKfLyCu78DtUnLzKtF3LxoVY1N45/bOjTSOTDowiXAJK2oDYMbRnwQBAaFWAO
5zp/b19p34nWGl/PmcIWlkZgD8MmbYhoqFa9/Pw1VUJjPAmAy2p64MxwJHL/4x0e
BviyX5EKKmJKZxAR4/qBVshyKA7w06ZROucYoOWCy416J9n0VJ4zRjAJDpgEHFsN
V48f31t+JFeUXzezOaK6BXhR/XLbHgejhQAJeL8DCeezo4jC+se1gL+C1/Dl9j0o
NxJ/CDqreaDnHbO8LQkdVC42RD+RYyRl3GM754n550EWfdpifOUoZqNEtvZmCHrT
qyLh/RfYjRRkjV4R53mT3oq77M+fvgTeBwaW478McUSVrtuHrA5F1oJsXVvtnhUk
ClBEmNkcLBaStspIIMdlwm3yGBMtPIiSf3TrhmxcehN19qgfP7qz14a5iV9AC6+G
B1x5Z2GdinKej5K/5aGsDQmy5Vd2idqOw4w5TEtzedDvCdGqRlbhRTKToxL8g9uf
iceH1xZRe3ZU1rQcW2u8HJ3oB6wn/Gvvu06zAnZaDflqLk6R/mcj7FGMxZh5vWTi
qCTAXfHcP4TB1TnQCRAYPRK1YiN+JzGtiXVVKCcRv6Qg8tBC04CGD8LV8wkXoW1c
bSrZbTtSW3zzUp3gSANTwabOtiNeV99/HYRB5ZgsxG+j+Cs+cQX+fWTaYifZGIfS
OpnlrDWKBU43mitl2YcH7BRkdkoCecVi7Hx8FcEZ3VpgUkOBVHl9sRoUwjGAp+bD
hIjnW/Y9VVTjXftB7XYa7oli4994CW82ffcuOPSvESU+Ux4w3FqRQfI195pV3nGk
P1fx8RtJ70ePKnNLH7zUL3ZERwg3QDlfiEQi4Sg4TNZNwXasExq8SXr0meCLH0pL
EmJKMZvw6wjAkwXQgC9n/hNvOlSq9Rn0YSu59mclC2qBe8gtjOAuUW38O3g3tZHd
30MU+hzJ/P8tgkoFiWcYbwMrzTNLA47s8pnRSl+kfG4spRhlYJlsh9x+5akhLruR
jP9A36uj/XIGkkLvOvAA40uPCzg46BundHWDbIl6Uee3ZWu0QyuqJIOwOgWo3XIc
rk0PcrvT8wurXipQaja3LFhsBGkhQrE6hHkgsdWNkGAbx1BzhqSlwJFcxv/QyptG
qlvXdyUjUev782GDGCaFWKoZ8unDSHI3Xfs66Wm74DBJj8LBcd8VZouGC77jaILG
hxIgl0Kuh5rWavbHP3WyAAafVJxjHOCmaMFxuNH/FFZojHq/8iL4gNBp1gGgP/Xy
DVDOVndEcT4eG/MDHomXoAQSBso/VVGDDOYLLr4WgasiVIlUbrQMGcWo/SUiCvHt
Sqjj+RhowUBZaZ2PCCNXVyB1fs3PLesXTanYZKUAmYRUDWyvn9DF38inox110flx
o93Qsir25Jol8/QcUB/h+Dhw7FqxCt/I1LMID7UQWY1nro0BsfnJ+xb4p7uTPTmd
93sP2TCTFuCHB6Z5zIvosHO7iZk5sR+fHaj54ffm9eaa6viDnPrS5kGlc+oJFrc7
HExBbsJo1HfrmTjQCFxM8qtH4VJXED1G+FXxcrzhjyuekJU5ZsnMFZvTO6DyT7Q9
bRg6edQH+6vounlEZabBAa/m5UC1QM4TvCv2RYig2Th3AL0kir5PxH9UZWUZn9oH
zZ3tRfU5E68z/CLuTjn+gVg4TzJipi0yJnfNAJf3+2/yr4qa5cEpXtpMUs6UJ/i2
ln/jMs1XH/SuFEX0Ac+wqU2RgRifUL/FKl02otUmm2EmCELic+qjrAesltFet3Dm
Lnda7kZxz1PTMXretKcTUKKFuN3xMTDEUpw2zPBB11goaKEtaRKbSDp8X0+ixy7D
HFU/VrrEoQqa6UzVXtD+z2IxToUC1lJCcWp0ZZS8aC34n3wXNrDJihEF2s1TWokY
iDtrOrLpr/7cnhUXikJXBPE1UwnXpigYyCEukJUFtg5Jxfl8kt4a8OyFF19tzGvB
NE/DeH7IqC8rXIaOyhQOP0WBpqV9dFpbV7YP5JS/ELYSXJv6tMeu7KuuAD69PpAA
nUvNBzOGo7E+SWIjf6Hfjs7CESBRuFw88s2Tm+KJTKnA8UIgmF8dakMueoAulHZ1
FyPxSJOLm10RvRedk7iteQ43om89+yqqDe6sxghjPzla9SA4AmP+pvrlQqBX9qrj
mOx1u0ZTHWMtRYkjIIvVqnTRvku9wsG+sByqJ7Tmv2hSkG5mO7i8CG8tvL0BDQYu
3BTe5SoFFXWzbkbwdDWwEpKHsBd5UXxOZf8Jva/ZFM6rzOoubV+Ceyf7WXJBaF2O
3JPyZF6EDdNiaDUHLalduK7TfIw3A+lCSwBTUneldNT2CXTTApNG4l1KGqlQxfJI
SdRPYw/78vQRtL3fCRxJEWSLeXPELrRPRjbNvF1NTDQIGslfY//MOfoXS5XW0WZy
4VAFPrI//F7VJckkR/iNItNOVAZEPjDOwX36Y8GnWClfO3mskhrDdxUG7ixOLxok
xZ8lAuQ6qA1AiMm/Dg3YBR8Mo0AyZovuXviQ+fwfTHMkCFHiQz/OfoPxbTg3Wus+
C6i8thJqTmi8prmi+kqhYEbszTXgPoI3oTfDd5BhienpsxsTPQqmPFk9nzysxpKF
HXiM/evVXSniMrgjHeNZBIy8IEc+iu1LDaJ2wdwqGGdFiSqCKD1i5pKZlFU5Z2aS
UWIqgr9Rc4czsMsIPumwivaxjIxVRYDeDfEXfQItquFvIKoEhBA8Vdr/kv6PyjnK
Ce28sMzfBeeXoZGaVborwNumPRU6mQobdSpP8f32c9AQ0KK00/bH4KTu3pV3fw+X
QLOj+AkymekXlE6OPOGbieSsQMaAISX5s4mDDTp0WuJV+Sq6eu/nIL/RqZ9lyxsw
Fd+okoFd7AA3AZC3bZsoNOCWAOr076ENgZ4f7uaHnjayGd1eKAIrech7uOcgxU3f
+gX/Kk25JgoyHy1hXgbxZIMZ249IVg1v38M96C9RMmqwxLQPDScmDsp8n1Ch298o
VBt3ajyB61zMBIsvMOdNGP/G5GAqJIqlxTcIRVV07dJ9c8xv2PWW25cM1BGtIj5u
obmOv4uZUqEfOe2C5EmjKsTKND9B2wHy6Xp9ZNoKziDIRH+aFzQeeNPdQLoKF7nc
bHTm5SN8XSTJyBP5sH350U+WrGosIbJoc2CVatwONM/CjrnZaZtC2HbDwNk2rDKJ
+mqZq2yeTJWWg5vk7wkl5I5AbOZsFqIUh3bVaB+OME9Rsevm6nuSSXINbHdp30Le
wjbVGJE1HxaeRCJS0EqHr4Y1HR+qFXfogGazvvW7HsFAZJoigIJ10AxgxfVxweGG
H5tsfnKdBmtDl2QdrI3x/JxRrvX6V/mTX3DL+6AaFleqip2IjcEDr52y9zxwmPb/
fReAqmEyWK6z7dWmlv660IMlEzI/Ulu1GRhwGQ37/u3jAQj2jCjlxFr2yjIQFgKP
gJrBDFJA6c/5KeXcgpFtWhkeLw/J2VtHdGFF6WBY+H0dKjIbeCV3fIpPKJPAsctT
99fi+ad151xADFK7iImR3fKkICradScVMjh2UVoKeQb2ct12cjsdJbb7kB+3HT8U
OFrmX6PtKk0DNPetiIeKRj78b9AI6cyYw4BK47svGLPqT9fEOSfC3BHXSN5p6I4N
AILDxSoGrH41ZUQg8CW2KG22/8/Key0iYyfqJgKcD7BeaBGBaduBsKWvaxyw95vL
bbeD6egSTlcHZVVgGbB7gqHYoRjoirNjLC6mNMMIm37gLDHA0DzQUJ2ZcZ55dzle
cmXjlHznmrYY6+H/v3Xz8szm5NBxYFyJ+Sn/1YIqYQmBjhtu5mZuHRa5WTRT13pH
B9v+BoSDkgixkZADRtD0Yvb/8vpcmCLpKu49Ww+Dbzq0I0YiK2ONc3jLFsVepJiK
C3QqxWxcAYXoKOo/91+pHvQtEjI/WwSh3eUKaMOlhHM8qej35TYgAg+j25ms/ylQ
++3APgG7z/+Ze/2rLTl7WT1oilrC08U4ApeFwGNlLLYeLPIwJBVFMW4JnU8bFBA4
BFYgrUihAg63VgIZ5eokVDXguBDdemYgvs1cN8c0bW8TYoGxmQ2WZjZb1NUA+dwb
LCmuMtS+8DbLCuOqqLkZtDjTJZHb4zNKpg99ndmRwURmZTEPlh8bU5LbKB+xcBkl
PTtrRc2KFe5l0eGBLUFPBH0PTbBxLdb0JXBt5U7iTWBXLSGKwn+2rBucuCQRGcHI
09OgnSdqQPPi7ekSYoD/G8t0MXnna8zPqvG9xeUEYhBWh/jQ2k24/1wqc4Bvhet/
IG/fsThvIT7oBili5D/d4CfVP15YYWXVAdyoUiEqfNH16YjGYl+4nOYszsWPyxyY
jP1xkR4pa6bGX+/zymw1sv1WFE9gfhsiQHaEJTO9KYGbBjdA555dWPueO68dJtv8
Wi3m1fvY5uotikrbavNvREl5W6czei2x/Z+clh/VIYc6ieh93M3sN/73jcL+xKTm
KkpulUUnl5HFPwsZV+43cr//IejKHI8XgxgBm3SHdQ16bMr/q8OVT4ouWu68SbtN
EhAY4TlXO36xmCoeb9ZZveD2dnlvoPmgwGVpOCjQul7zSctpolAajsxfLhJV5MMq
Z4GXlJYvzzn5zsvA2Mt8TxyH+JhTZ1OGEdLgtrOt47Yw9QhVIHAT8N7K9j3TSjIA
VmxwtCikz0VTU8XHnNNedTfDZYdtns4Fgbu+WCvwKtXRPJ8+5z+LqOC4S/+gs3DU
beB1mCP7KyiiydoDJeFKWUNuPForm9qFVY2z9wD3MJnNycOg83cmzF9p/ZFHvERV
Q53D0C99SJadaXNjQMalouv5+PNX5XhhWecMWDxpJOHqXF8urEG5XekUegQxVhkK
t4QcQSnwqmlqpYloMzULZklZiNyFEziuYiew49cYWH1gxZw8szawT1uMdo+LxeSe
GMEKjBTBR1gWNibUmDAAEQgfjjEZ1LKmhUCIgpmuWQPUr81KyP8yxMSLh97AMtD9
md9rg534rSKrUgsUJAyu135ShSO5aSMFPqr49qNV7E1hjPbIjwsLgDrNp+tPQnuv
fJORZVFmoCA/jUGrnOaQiUiISBxQEPrpjpGX6uwtivMaS0LHytNJfP4LUob5PwS1
QFYeNoIMrzsuBeew26QigKM4y5A0CSSwBfijuMOrC47sQ85l+rg3Z4/aZpb5W1uR
nS6lkgTW6VVZISMNZT0gMxhqI+riOOKyuBnxdiVKrfzCzRWwkZtIEjOBgNzjgFXM
GZbDqL3HQTr7CPlsiienIxjjYwJEB9TVSYFCeDsikDQ49ca0momFNBqimBJ0W/hP
xyVsE9kwH1yDmudBdJkCNvnjSNSCSugDxsnLO+4s/JpyFkmXgbjxFHmSIjMJokc5
cWhFS0/GLzi9vL7xI0AreRuUClm64PnYHmAamBevL65K2v95LJ0g9exiX/TIbSiA
YIAFbCbUUkdE+Yx1xakQop4AmQr7K86IFqQSLkaKEXgFPN7rJTNDkkrmzIozh8ok
H3jaxgNSh0t4RyXLkeseTikdtJIxo2W5doYU57EG2aXmTeeVGMrYS2U+nww6wJOP
2sZAlC4zhbE9kNM9TDMpYCtYtOZEnRS+0ohhOZzmEbTFr7sAShA7CVS5Rdf8U/TZ
P7buBzHYjAx5KpE+w2d375Do3V2OjWQygbQUhWDGyWmqeIfGMktNgpwj+dxhsznQ
emNy4juBND3/ih4Bj0iahzgxOVU3wYVU2wF2D7sOPDx/sFI2hh1pzS2lIYfAhUwG
/dwr78xo42GC/WhgutvSqstVuQGCEX1+6Luv6l32L1sHjm7pGsS6+Mt1tACfbZF5
wpqI+StgHnCn1q1Ng5qPIZg8BovfLXupxW7pW7fFXbNHkiuHH654eytKQ8Pzws3t
ZBL2dK0Kplmw+pYRgjMQ+FBwjeBqb5uIYQOlRCD/N2+R71gu6pROk240DtSlO3Ws
XD0uxSkWcznp5IL/oahhAM5FRgBOA6o32i82CRKXXACv2WV/ttvCSPlleulgHhDY
65MT9jD2Wel9y3T4a9gF68bSkZw/59UD0ddiLlbsuEjLz7ZQDgIf3MT+UC9B3M5s
vBM4OBrXX+Qzfk/FOFTGg02VOl7tlmq1ArqNFDp5kIYafcUWZIhRCXmgmOc/WObv
KkmN+mhoyGbKJwAwUBWhygYeXTCLZrbE5ZT1wsrWhZufa3BwagzKTrjJdkSRzZ0h
TG9LuZc9t7JEX/6VTo82zW5+oN1XAb/ydGHIR+OgNwWc8wjfTQRusft2F87A3Oc5
5cfHsuz6UmWdJZiraczaI0jpBHJA7lxQpaw9F/Ymc2kpMvB+f3H82iXB95VdKYYp
+bQQmeWmLIQRHyMshSmXm8d9yLVzMBYcPAPv4UzVxUI4/CNKIECHvB3UG546vnDF
9+PUlEMExHQwJsvYeXQ64P09Puoiy0mCTt0G54AlzbbCYrEW2kitAoaMuQPHLlrM
y7j2PB8uExwcDhpK+hGHh2jM+L5W80VARJUq96GkQcDalvoxDvV4gddJsfubHRQe
3KhVUPd/GxPrSlcELWTg7Izi4rQ6JnBdBa9URxiR2/7QZpa1dx3iDler8k+pFth8
icpWoIvW/AgH85z5MitAQlU96a1myI5OArspc5VPgOR3AWpbwQHndthXunwYcZiQ
Cq4YLUIwk3VoB8JEyz7sNdtamSdI3p1vqY50+3xmu1rDnBmz5qwhwEx6ZmIHl7gN
cGwYgXYLmsAJUEfJJDoo22tPKPRCPZbRje59oglbk4wFUK1BrFs6NmA+v/jODOPW
VKDH9s6GzVqzUH5IiJKKjswHUmDMr3O6jUqaA2qrcxucRHB1hfw8/I+q9zTDsjCW
LE0hTyzWlSuWBwV0uXmG3FkRqdDQtts+E5pckVLK5zjrnY90uK6Oy2eVfSwW1BJO
dBBPQJ6YNp3vWSWukv/y/Fh09qC4XEE1otJRE3f9CVJOD34MJOAMXk125RzadsRy
VWicaQCj4FM/jIS/8kWdFIha/q5RaUX5cLuGAJuSbUGOAj92rNXYUo5xHcU8qi/I
FajSG1f4U52UezrEJRbJn/m81xZazJHDMoQKE7DkxEEUAkTt5FzXHf73tDpeW+sf
Yp+RDUx66c/f/je/CitmLNyHb596FVNF67HqsKyhB69CWP59MUfSEC52QQQZDTV6
T1i9RG8Yw8xIPsCilfQtCb6jU3sISy5EV/Cmq6LYKH/2ICN46mpHVFqdGRWsfOT9
ciY4rX5F120r4+6mtAzFdn+XxFlTJ2O5avhmBMyjRcQOU3csq8fplN54am6wy5aq
jB0IFiJoUO2ukkHY+f0l9z2V2tISF16hqUsi17ARyLBzijrDSKry+P65XocBii8v
ABFBxobdoqbYkYI8N4r1C2Sc/Esu+ggXBGrhwB4Jd75IWm8RKHkAL+5HHRekPCj8
wJNfrrvrS8FebXzGk4oRlwEvl+IOenK+kSqAYumv7/YDkufHGJT1tfbFDQO95ktP
C6kcCd7HNd74Kr9nP+w96S0MTsUd95aESU8PUmwlIJP4BS1x/7KVhMJnBXHr/c2q
MRo5UM9kjMGxzB64COufUO8cQnnAb20bCf/3aJpTAcyPiHkE5pZ8oop6m2sol1iV
ihsDf9TiV0Jo5YNO+NvNDgZwy7psbSZgsoHAE2FnjYFHaDGuy4kI5sVenDrBV3LF
Abtn1t1UPxUB0Vc4+sDfSOmtLLlNaFkl6v+PXou9Qw2qqH5K+3HOUu87eAA9nWTR
8CW3VuIGYFTdJWKqVo4hj8PpMiLwMtIR16qB5LZL2OISKALctcoN9YeD/MHDi39j
GZdZazTzQU0k+tlr7pQlCNugKMcTk8ApmB0BjtvWeoK8MHP/XHjHcZw2KVnNvtfp
4dhAp8b4I2P7FyKYUctPbemikeFUmzZzZ6sFpfYihMhYNkBZYM0LrSCYN53z54Vr
kEGsedFMc4RTbj5ew2e+gAa0IXxsA1S2VqgA8DUNFE3DY1EKbQOt2E9gzNCEnEIG
F/6wEYY60W5y/pTT6klL/jIm+SxjqHY9yrYZ/sUzHAIWIu4deFENiowqkdSpg7e7
7VkZY2E0TDvirZkKw+Ke6Y5I3ONh7mR5C4xXqoCt/aVdAZS4ui+5+fQHkG17fogQ
QVky7DQaMNtr0qazKV/r60FlXBZdQGl20SRCUEryxIWsa4HB8Nj5/NSiJrkhnYfQ
nTEt2mus1WSgBTY8G4U8qrZPy8wdJUMJ/BPk6KUPNinNVglsBCw8ENLF9JfEP4qK
HziLWgObZBAf4rosRHYV8r5PLxJolh9zS/dBvwtoTPdYtJA4Y4ISduVE7urVVYRX
jwcDxbaDZYVM4XnQHafDFwEOed0T5wyY1eE+jvV2ejd5IH50uPorcxVQ1k2m4p1p
mUEE6TbrbU5AONXbaW1fCP2BLvf1PEKNFVP2YSYRWejMrzMoj1qnBc0yc7gTPcYk
JiwNg5LVI1hFQVgMvin5XgWbEwRYtYZV7xJ0meilKmUkGgOV+iJ0Lji6YQe3x0Ao
UG5b/yIdqX9TVI20zfrVfB+KSwKoocccb8Es3eQClzVFY9PdnQF5/e7zoxc9zxOk
dcMWsIwJroIEeTetsckILQ9Wn4TifA7uQxPexMMTv3dRnT+cIW66c0ERdyCT9aVO
FvJNvPE7afutX+33+vCIkaeuQxUi36TgrFKubursJL8nFaqv2WkCCtVUHdgjpeCr
6Llef06C6fuJOYmcha77nZLRHXr6dQtjDmpfoYvPzwEmwFB2+DvYfky+Qkvvh97N
mwfWcDon7Tmqo2QDqt/vbFpG52OBcH+7gwqpF0S4jbluIc4+RWkhScqOJmBBBzuT
/pTvXY4/HgR+6Nn9KLHCPtKNx+A7+UJsbgTYN7VEwAv/biDtZLEMZ1azewZUKJ76
X5/uJB1u42O/2FuaabrWaaVPhyfQe0U+qi5CXgxTLjCjWz3LzNAjZhW10BCbD8W/
cx0oAR1hIbti3BMciwP1JIgxF58K6QCBuv1ih5gN6y+uGUTZi97wmmFaGqV4uggs
8+s1EnIsGoXBCWUgNbjYLDMHcETtY+kaEIgsXBJtd8K3was4jfO+gvR/66tmrwDr
FBfgj9aWs531RdAVVFSZei9TUWn04BUX596EsArk2l0hNDJ17FdMl63kM3uwd78+
/pTN17ysNK7ouoKsMiKbY/FnV/CVReItKJrxP25Nceja8L81DQLemX9524pp0YpT
BGrg/alDlyxDRR2CKCnCMWR8YI7SzOIyXP8zz3T7kwD0VH14wQERs4rIZkLmZs5q
Lkjp2Qwzfl6iXmXx+T5x4R7F3a/B5P2pSb4rL9hh6xbuisUAQqyKlMM1RNnY1nmz
fRPA28Y2cSLBBCvy32n8vU0LucBtaHql9OO9dCH3FaAbQ58JWdtAM8PPTBh0TEek
riLm4oib2Am1uqwquE3FmkobDoJCtZj8yFhQG5M2uKiPL+Ywx28std+lt6MhBlC7
T21xo89SAoR0/uKxZuu+JEChdzYcHBiDpOOFLM6gh5aJrERgkrA39naYCyz0rAe2
KBXGX1pQS5llVAbh2DJFM5aiYDw2nxcGUahLQBAN1HU6J3EvnlyVo2YxaQ3K4AJF
fjNMnqEWnLL/xJCZJZKx1Xd3o4KebkgGQE7wICm3OU5ruQ+RcvW3rokEZOKkIgDq
9CQgiFeba1du0dc6ncYCNwThZFkvckxGJUedib6N57HfY1Ln1ULFKBEgZhwV5N48
B7gXmlbDEkNW30X7Y/G9mzktTnwdFrty2xJtP664QVszRZ2DUf1AYx5Q1ALHgG/6
xmxbnUHlXlm5Li0lzGSReV3yRdlWUMPScY2+uixCXPiywbG5WRLbMq+sYjAMy84l
9vVx2ElmpjmRfLUBYalCMgbc7JMmG38q7gY+YTcPkSEZaF7aJ8cRW2x2sTQBRX2g
xQ7qHDU3g9WWo1/7nbCvFyFZagyaJMghrvGyGHG0gbxMLJzU4SXuaQgQfMwFR+1H
WJy1dZ6vsutszQTbxAtTkLOyRjA5PkwRnSHqSC5lOBTAfJT+mlQ3BkKttEjD585Q
StoGaDjRJc0WsDoJM9QLxtmJf+6V8xzNZ/OeC+BHEvCuAb/awOBaYfeddO8u7iSO
gA2SAwAFtV4qpdGsBjtKcB9eh1PS2U2OxmaaslRqdKtGek7Dofb16/6UqDpWI1sR
7rN523v3T37SBHmM1EadMclNWqMWpLoaWiB4e6NUUodHaF4fMOESbiehrdOUznd1
pKXJdyM62YsAHVzORaHlIE5/6Me296kqRbo2SHdko1Z1G1/MAB9rwuFo/3WJFjmL
uwz/zWorD552OLKZN2fghE2PtQC/kRu5MB7QYMUwixK3InlRb2YwrHVvnfkq2deh
pFMCFQOz8Hu/qBEGEeLySup5TQm5MPVfcL6ex8pbp12dx1y/bNKsplMlOaU9O2bJ
H3d9sUAOD8gWRO+m/cDZCUKiBYinbUphXO9y1pvVsQtpOsom/bhLFPHegIcjDqv7
u7caE9mI/d74Dzew8aQ3ak9dC6b7Z7CJYmp1C9lIrvhzAPJrX7QV06gTSCDtwZhP
mBvWw8sUKRb0HlsCZD4AnH2PI+hbw6tIM35RZ9WJhL/UXIWk3x0NefyucLXsU4CQ
rpFJI1v2Z4+ASNa8A8EwfZYenCPf/04RVZyKG9aIGjfAax9u+1t7b98suwa5R8h/
tMMjsEdDbNB8YL+O9Ky+eAhIRfcZZdUDLeALkgmbLCTJWVDtDSozLST3js8PB6yY
992nWcYQ71lELe06dubTpbZRnJ9LPZrIjrJMdXweJhlRYnfqX8a7A/cC/ZAKNZbY
vR64CluJni8TJrDXo/iQRMEPwPf7UjnA5sPNGM3Rgd5hUk2kSFaxqHpmqBs7GkHQ
ekC0KCXRZI16DA5mTjsIffNpd4tKjx0+nOynRlB0wbSfQYIO5YBf7GKGeLVrlYBv
RMXGMxJWrNL1xf4BE5w+OBOdRcp5bENxwRYCuymU7wp84AADEcXvqikwgGK9cAyf
+gl369pnTIpBGzI94lvrKX9gFBfJSr2gEHKN51Nvt9lEwoRVRbJMpUu5XvtPiJxc
HFM9t2PmQRzUIA+zjR5YrFmuT2TdOfh+eJbajgnGkR/t/oUDFgg8+yqR0VD044De
pgx68iKcM9E316O3sMxOFydKY+TCy8rxA0Ws6+XVf4PopZjfHdxXGnoqQfRfYeJW
aa2i4hA1kk/meYoFQDIepy0YM9aRUpOFYCFUsrThoSunu1UsJJj7t20t/5oloy11
stvp4CBNAoDgr/UWfz+naSfEfEfGLuZNpzqRZJuFJewix5lXXqGBts8r3aHYe/PA
e5TTv1ESLnzAWIFpvpeZEwxmT4NFatOtIufOGP+nIh6lB3V2IWAmcnVQgjq4oOqL
SiBHms52m/1paEvctJLVYREPu9NB1/WryUnQ9szAqoDbnWWMFCIRcSF9gqT7xFI0
ybKLs/VLnF4t6bokIRKO1Hd+dSH9QNgc8RnzAJkK2y54a40ppqZp5CnI2YhXB3By
OH9huGDNzoDFIv4F6c0kejOM5cESQQtzUEqUlXCaIp8F+Rz3vKSqE6hT9cSE2mZp
Aije72/ztTwL6czbyE+tOHxWhWe2MfHlRjEEwONYeDXZw55+pUs3r7qV1cULd+DN
CmJpqMBKoYw7T2s5aQnDZBuA+GawgrfbNvWhcK8b0NUY14erqLbLgikIVsdS8Oqp
mFu/V14LiIK77Uyc5FkGnByNhjy0QmXBNTwy19JdJuZlhue7Hi6Sm1IdZ65HiwSm
Ac1fA+ffInIVr+yaW3heFqJYJduUq1EKlJPPJDiNMeoh+V2Jol1tY+fuHQToO2Pf
kPogdLHJOq3gXuyohMMMerMTQ0JqHGkT7pvw8VGX1dXWmIlVm45dnTjQ9+s58jtK
W2/7K2hrO7jaibQ3Zsc3sMZevhUphPwdC+txcSLmopDRqmYjuGiRNbOmZJMyjiua
/15JQME5y2ET1yVV0S8JEkEq6W6zWKQYGQXl5cC0kqlqVG+8jzskDfIvwwqQ9ZrB
TuMw9cZ+npGSIzskkSsztqaHa9lFlZvah8+p5i3EwvC/g0Vq4WLnlfTViXxQgjzi
/PtSWEQzSCHB3WD8jfFnPY+duABIxAObgfLhQcNVVJy8AtPrOAKqvbiF9KrXBONw
f88f9hvt1tWJUvNtpSnQYeBeiUok19fl55j/1SXjPZ3ld7H4A38gTmEBp/w19ytf
LMPu3+tf01ZvwfRA/c1cmJ/Jk6T1uUnwWYgRA0nvcX6AngDlKKvvDW7WZfvu3K2n
Xe1otzPANHpNHt/M+DCuXXPwajbaVn/UD76zew8+OgIebO4mOaCA51USE0CYfC7g
8CWMglFDa6JdljhZGaSyG4U2I7Hgr51cgAUQUeHMjYslvaqL1FShQgQtIosiZ7+9
x+8bPD1qeDObaadaf9N6AK+VPKb96ME1ZtX0BTYKzm5/PoHHTr1XUWf0dNJE2puQ
6O8oPho6QDEXkIUUhZ1WwcND/v02gePhtRmJfCaXH7DSpN17Tkjba7thljDQwS2J
KPiuz6ETGIvPdWmuiQlRsIo5ey11ODxjLFdZz2EhFkamt9Y6+Gfyo1BI3KB2NTM7
PBMt/Thlyodfr/jWwS2YmwjKyzIeUcWw/XgkeBAbhcjIZcJi+ndQd53pif721T/O
f/+mn6VI6+N55HfcBJZbN88PZAkhJOhIpK4No/FuSdWpUkNouxMi6bSf1bbuiTTL
OpOem0jXfNya2HvycsQSjjZTX1lT8kLfLzf1gF+4txMHev3YWuDSIW1Yy2ubUqCQ
jqHR6fVuw4Z583Pl/fUSuM1tBXEg9Fluoi1HJKrCuhN8iWMdogg9zqcIkhK1/ttZ
TFgPWqjTPJqhSfSCI6tkWZx2f2eTjjN5MBcfMCTYoN0BwILYByVP3dExMiujNIoC
2kABI0uFTj6YiHnF25YDTvORWSFxDyM8nT60RwIx3ml20TPv8lwhtgVIVh/mr6Z5
78ha/llTWNpoAkK68R6Q4hMivjq8LJ+lbdjfaTuSIEk5sWJxYqpsEZzPPDma6eBI
w2i1gicdGkokrr2L7Z14lYgV39w+Pd1Uve7C8exdh5yTZKRKLcAYrhPzJ3phPFbb
RtTAkYVnaKKT36Xn+G7yqosQ9we4YiAnS/En/yWM/+YMaTBBD1Sr31Sc+tcv6d5/
0souejAv7zFBqowJS9nrUIDZ+8CLBp+6lN+LKSHb1FVt276m92IMUIejcp390ghj
dEn/gdq83OMI501yYQQbEI2x19e7YpNLwo1JaaGJ0pK2F5Wxq5IWH3hIo3ZGggRn
sOpaMH2cAxQj8lbeNYZOlNyd/VxOHTiK2rtlp2JktaLwqVACy/O/9mqbBbsJE7fi
EMGl6HhRkMY8VmPY0Tx2msvmC8nSSOCodtA5YknJVIzaBAQWX1Ky0iMAWO3WqmJd
JV1njrpcvDhnhClVlVfShHef3LZwK73zWj7MTDXPIStOk6TFE1YKSDZz+njmFiRY
Fkb6Yrd0dORZie0Y2fYwkLQzZ+n5rzkrh1OdeBz+Tz0kHJrX9ru25C5koSBPf9yO
r7FtjnUcsHsVhX9hJj4IsbYR8h55Xpcl+mJpo/kOzaN2h7IcxZ3EfOIycbi0R+N/
ZrkNMqmN63l4z7p6yBRuN1WhaDddMQ3MOYSEGFpIs74RBcP92oQStyerf23xmuR7
wN/SaAdi6vbRg9eIZWOcHbBs7GwuBIG9gPInhCcBZ5AW50lBB0dLgetcpBnC+FV2
/fVYBeX1G4Rvgyt/lOsPCPHEU7XDwpTWxoWxaLrjg+kq8MxGkEOF3cD8Nm/GI8JF
QgQxkjSTrvvdnwE7ygxKTO8VLOkLlHjfHG/uy7RXIef4xKWckTOqyVjdaVUDo5n1
xndrzNfwN96UlR0XYJ733hahrWHnCoF+myrFJ0oegpUqASXqbUu8qKGlWB5q4ylH
/mgeS1/RG7jNy8az10E9CDN5/E1gYSE2uchyVJijg4gOpU6J7hOq+xYFOo9Yx/U3
aOrtaXOYdI+5L7+BdbkzGIG6uZstUnvfvnBl2MJ9wrNMCvp2XXZBbCq08vU3hOKh
3ssoC1ClKTCwYNV3Rgrj8xir2oSSEd+NYIWTybi3pfoOBmxjSvE0WUI7t+5xC8l9
czJhWL7a1MioqeAHhnadyAUAqb7TEZT9Wcfw1uxX9M7GJ4zHqrqg6B8AwPGiOQXx
3M4nAWsd4QLvVpJAEJ6H6azZhjkWpJtG9GVl55Bkb33MOsmAhP0vVPmIwHoOMmv5
/In27k/UGrpTf0oSeYnZvrqGYCehn+nR88C5wX7Kr/+m2Mf4WylHd9xC4b8RImbC
RKUpfs8zlP9/JfT8FlStVSOakMb2h1NCk8iA2pEMcYva+YwJwh7qWe08PNVaWAQ0
gCRfQfO7a8tEJGg7WblWWerohRxzzcsjUy/+7H6Njs5b5aS3/vtKagQtL37JdBO0
pJumSH/0sC2mw5geO+qjjuxI7EsTLxq5sJNXqg0JRjgjtcHQuYwFQqqzN8dHY+xv
cMjPOLZFx/9batXswoPEXu3tj5x9VqwQVTopx5n3F7fWc/K16aPpdBYbAWKcfDRg
NM6faJ6Pw74YZnMdvpzAlDzpD1/kfU2SX5s5Z0ohZEO6wy9x+ARqCYmDkD0z2+hV
nFpDLv/5Zf0/ZfhH3sdkVA0w+HQbpUNVmNMDTrOAnOzml0yTze2KQctdKOfJ7qAH
QHhJaTzKQRPzVh8alVufvYlG94rCrqoiPCeYjIy18ofl/nTntVHan8TmJvassirt
KZvl0494yEzKq4LjmLzzprZyF+dpX+q+9pPkJDD4lvv2eb2qtCMFpwFcpCNoG42v
wqvrH+Wf7nbn0pqB1JnVvyPymTuSLOGS2I9k0TjJJVGQli70T04yD/bwmyt+R9vD
HpFRDKKaMVtswWJ3j69jzCCGPbHjzn5M9Zgk3iUS3rWeJW2rDoMq0sYV++ByfMSD
3mFeJh0q+jSc0RTgeHZ182U6gHNB066MMf65zdoqrmpdAfxw73OfjjN8T7ktZpy0
PyeO5Kphl7sEI50hxSNTGifMab0sOBMh4dxJcZOZOqHFTHe3G+Js8wqUDFel7xz2
BcXx2zZoJkD/hCgXNYh6Kyskuh+pyLCvLuXihf3oWKRDvEOr42BFr3z++79jAhvW
0W+xFeQ+j/yuuANLdsLTvMk+uZ+8E3DqSfhuzb3umQfBOqblap8vgI8cqVLFXi7b
VSy0FObfxrr2qw7hyHhfcymqhfXIjyhcvbWsgLHg7sgrHJfcpfroEyieglhBLIYS
i5uEnBEnLev1zLo3yUbfQNEG7USaJ9gDl4MV//aC/F+g0xlMrZe/YppgtlJQUHKm
y0ftTUBB9XmKO0kQ7uPx0EbNy6oQ2DuEeCb1NG+8jYjsdJCM36ZUoRLJHFAtzwQY
HMcGeRkUVg0nYIg72GpSb1/zvBrOQM99xnPnajqUYSZglCMySR7WMEYxHYH+/+ZU
c73odjDZ1uE7qsZEwZgTtDhNDGa2sQ/KOnTUVxjHSCSGramg2PBUct3JRAx723ER
UorBSBgPy+8paru7/ABYBh7xdGcLdzkc4UI8urUXO9M4dQ10Ez8sK53CjvxOFtV5
6FgAu387jWZZKlOEbR0VtoncMn++ZXUVf+LwtKrxsfVEXg5kvO+Q1sdt5+hXJnc/
3OIKfWDiIwCo6SPFEpfDlab6IlOh3SmXRth7M5B1lUpKjJNkrBV4Qb9QgJyram7U
g60RlfTHmkKdeR9GQSELxytWXlR91njse6W2tyZ6AKDdIqbRP67zuFeRB7FmHzll
mJndu9JVSLQOnopmyIl+t6Bwgr0desZ01RlQlGw70bkeBD+QLDjSgu1dKZZpel1q
pxO3kNR+ExKpns0jvPtI4/hPILHDByxaCPDfZwW2hizRtqalpvKI+ywkuISgoDyZ
QqDXR9DKHIYGQiFLJ34CGxvgHbjGaa1kjmW+jPpdWRhwf2iI/ld6gB9VLjEkIYl0
V7uCbS0saG5gfVmijoGravzWEqSz4YgK/21eVSveJBD51kpS9uU6Bcj63FJb0t3H
ouq0RyMgHnJhUnyKxITA6Eg2um+m0VNYehR60YlqscAM3jtIauj05YISyZD6IZ0Q
BE4SDjwRHKJc9+XMyI4mDwpgfuPRxvh0oK9WQhH4WXyv9DryRzA5Ty0jUBlIvJJ0
PnDn7O6tGJCzf0qCWk6DXQgVbgcBhwGq/fcnmpgMjrFP6/apS6NqpqMVZdVQU5Y2
p17yJ+BwHZ6KKAUt9yRuh/lymYoLZg8tCnuNhyb0ZQ3wh0jnx9CKHeLqw5NAdE9C
0zurikefzmOkRxV+fSX7pQvVUOJmzw2HwsKKPkNnCPf025ZZCZwOIEWexqwoNkxb
OyB11pe3qI7napUECX0+3icmyTqXycU5OgrfiIshb4id/v1alxyZIPNCGT3jUr03
dvk3jOnUUIAy3nkT3SJJ51Fbs+DosFQcj7xoQX2orEc1aw0C5/cjJZUv8E3Rq6Lr
+dBsuYS0fsmFjfnShULePh1AXXV7sRpmpkJvS6u8ja3anXGLRT1jdvy39au6E9Tx
v0eiiDoZQ9j1eoVoarsoSWOz/iJ0tONpqRjnnpW1EJHGhfrj+yiJe/iBgu5NrKcU
xFOOl6ivbGGzlko/CpXR3rkxrpkqWJIoR6LMMtea+xRL8BCqn4g+nvVrFNznZrzk
BxjPHNkLdjpqzswbEtteGM9m0VFkuodTTtqzT5dGuHymY8un2NWot5QLfGYNhNO1
/xTWLCVPqCm78wdI+cf3dUxI6upLi3jjm3DAbzecmzs7hmgedcbUSC48vPUUU1Sl
am9j7LU8OJ3LxkRq7yAkmJ0ZWL0/x7TMB4sX8bFMgzDLo7hH20pH1Xa+qRhBDWQb
E2WT7MWxuU56BfdlQwa2GdvJwcGZxGc1Q0z1fN9mEhhdlsqDNsBsN7EeLDqbjbad
uKHe/H8KdS09XKo2JhyZa6j3oWTkI0anYaJ1hKiWZjQu/qR6akhfeMYp0/dbosgQ
K79io/Z455YlMwsAREUIcIEeCWPWtXjSBMwhlEUOqhXpPyJUfuK2Goi+PsX2+vnU
aT1+p88FT1xQoDqS3csXtJ9Mt30EJm/QKhBkqKy2TaIGNphgXC7OkqK2kAJL6SJ/
+/M9Q4Bh1rrAc3QeO7K5ayOYoeySpzjQqaOT20rbY+OFkP1M1+TroG0aNxVMDqqH
OzE95kHaFsWqeYNbnnsRT148xtJUv3YvPD13K4I1EIVMagdKhv8sr9PNgLgsEoC2
yYPKn1FXgYFroCUFIaMHGNvgAUFzwXG0mb0L406rps7Jxkqgvb5zNEOiZGQS4bcl
RwCmuoAzmvKs5mIn8rHNsIQH5ZL+SMzrYyTeYTkmQwtBHczMJlzldiyiXqISbkZR
IyAenJQfyWkwvotqj9DVgeuxEKXGsnFtUVHSSUlEISvp3XqI/53C7K5mkED2JT4n
XMLTt34EWmerTtNKpYMF3Le2AtA/kz2Cg5+JiQUTbHb6mbSSZ3E92tmxX6rHFj6e
R7gPAmK/0y6axMXtJuY9jXyYuFchp5pkzeE8+h0vJiK7/7gsL784lb/4niYU2KCP
a6+oBLPy3KWlQHsUf3V/FQ/5fNI4Jb/4Ed8QpAUc64Tx6ImYxxfgqWwVa7xPaGj8
3HuK21why6JkQKoC7gk1n9bILYuhkr71FBGifpZ4GaVK37vV62IOA54IVrVmC3QF
XT0d1Tr/NDRNQgbHngZjOXJ8tL1fmfvINWpsWVrMeVC9zHZkDnbHDiJT99bYAD69
ND8T29CZ/Yyxduyw7QzR0QZx7ET7mAy2YRsr2svhbDveaJ9h9pURzeMxYfbaEYkA
RZr18lBTVx949v4lQkqTpnRpWmP+g9f3WAhsHiQqHZfL0rnjbYhzqlAYUyO4ZvQ2
vo1zgmOVYeR8StdJXYnhNXSi4+qRZsHJqfRaghrWy0HCcZSKljWNTF3XWo8j2AFm
puhIw8XkBGU67G6wGqD4kP8aYT0VztdL9gCqus1XZy9bzShwc5RXULZLxqkMhtMU
t6bYuI065TNCXv9QmZ3TFQ9z0Um5q0A/Hz4sXj88eYGEhUZbEOaJJtK3pG6AhFPA
lcYfHTlz/sC9hBZOTYxYIHLxQyBWw1uc2MofTi60J3KI8iG8dpwubKTUWl0t1eSM
JYAOqrt+djeKBwXBXjJlkseyQ+62Fh7QepciB/xiPS43WOXjuwawqxZFcINvp1xX
7mBM9Jk9WH6oovfOhRVKmGj9zEFHMrjYZMF3d1oulirZzj9GPylgYi58vLuObe/r
77nEloEkAFFLGus9dRVbaKpgFhfvUkPK0mXSOMgtNsgNnWRNz5VKYTweKbBXTAGe
oBGxrsGhZzp8XVlSQ2zwIV5TUFk3eCvRUqyVbBwizrmnzVj46/hY8Y/zm5mcjo5y
7nC3UjEatWcKwhngrfLWaaRcC3fTNRbBzi+jWRu1UuCe8EDn6Hod4+j0O3fcP2m+
rwo+yjOnaNf17rf8/LbXrC/1avphVhVlrNf2unNRT9KJ+9eM5/LXxh0oCYo/mn3t
a+Z4l3dfySETESvChekkxINeRVY7HvKLZISvtuuGzuUxVCWU64PSPe77JqkxK+Wm
Au7YqCppITTLf/bMW5X2IqvlwBbgsJfIZSy/R8ZR16BylRswojAocYtjAZTScQxA
63KOibzYe5+KHyGGgSQuhDu5nqZS4O9Hj1MO31xvRnB21SzE5ZgC5MoAwHHrPiDL
UNhg+dXc6AJJ2lECoRhBLgV4egZIrq1FZUP4VeuMe/WfMiJQEROietdlm5CHxLi/
my9VNJqru+u8PnhfGSYH/2xPCxXHomcPROWDJZ3Qy7Lc7k1UCdMwh5lFT9tYanwS
wvil2LrKimxXwHsayfVshECu73d2GrlU9YdgklJPtRZYQDvqB5tntbhzCgnWJbi4
2r1AW7NDyX4PLp668znFB/zdA1Pu4Vxy/X3g8lR5WV7sLa0zs0dUUD5+rxOPC+zI
ODe/CVrdGXKEUge+1w83ideK+n/tDjI+U4FY8o7rnAeBo7Ahrr4MBHIPtUPBYO+l
BYjx7xa/TPcHd9FVhPuPyIW0iZSyMcYudHyQ4lXE4qJNTov51oN0nh+OL3o66mNY
tkGkN+Nv5ICRwLno+RBXMHCRRkTCP6oZUQELhcdRD0tW5HW8tp3669c3HTK8JFkG
5dEBHpyV/lr+CDqzdAsnzwxJXlhUNrtP2DTXF9wGl+Rx3mG7+/rvbWC4W0TNsEm9
fFnpz9z8xE3Yp1svs83ryBi2lk7GZTyR3FWQ9p2axZffZ7s0sX/icKBVj5Jz82xZ
zFEDuH/vaeKHXCHcVaP3OqXEe04tYkaBnYIkznqhUI4v6tFu+iVEaynAzzhO/eZm
YbA0T11os6BdxEHBeSg93V9SqU/htmKV7vv3X1nGihONYw6IadjzxGkvXwpxtEld
kLNuvBrBr5mB0sY/goq3kwlkZuC5/C9H+DgZBUYna0To+8EsIeoxdN99q7S/c5Jh
C5i4DRSRNAYx8vimpbBOypkIsatOuc6syL0car3tAylhRcucDe7IlewZ1lR9tLy0
/aMdOd9/Mgyq88YIK3/KF1m3KpiOldmV7dT0zXx9Ku3LLYrVMmJV6qMflQKObOn9
TUBZ4AUOYSD5u7RdLHHkEW57ZSIoTA1S3a8tT1VS3X66zaJJo0VcD5dMBFx88ZiG
cqGhNm+7nQLsNJBRDl+ZI9twNSFNUr9T+8DkmI04FOHzaeZtOYv/wfJ6y9g/R89+
QedjHUXc4S2T1H8QHOW5S8WqW7YBkiI5st/EQZKd0/Ju2eiyJ2JT7lXIpcAipu5D
6IWyllPgah1rf5UilWTWGOpScF4/vl5IBzsnMykvYt2q9XEi+835To9jgao5vYb+
H8gkipHGvyIPb3kmFNz7JH44f9hQywYPfIDAKzRUhxU/9SAYXtNi8CDMZdB2VHIm
2WEBr/G8QQvdyadqZh0/CY1qvG1PO2X2jjEIzTvHkks5tGv1j98ErGMwpvyoMoyX
3RtFRbP7ugqSzWOUsUO4vqD0l1aq5kV/3ebiMWLAtLigQ8Q6j7zMe9j/wy6qwRS/
A4RutJJ/a0c+5riaqv9EAddyzWXxTQ3WowJOyUv1lVFBO55JnEzlUqtNPL6ZECoq
OMrKYbkptfy2EZ/fj1T0dQuzFU9fXdbdMYtIimZPnKOMcPP7rXCABppPC5MZbhFR
wT1NeXbRcxXtRVMzuZNNIMymNCNjQaPWh11bq1Q9DdmCPXLB95F/96zmHvmFaRRr
ZYHetT3T4P2kMHiWvJvsrFrbKoec1sHqNMe80XZSW52f+Fgh1w6M68dGoPd1EI0u
iSKYqj86Q3XqIRuzvtGlJ9NLuCV71mijRkvAPEJOYpLnjSWAPXsU0Qlzpq66Fg5M
LSDRttuXFKP3p2UDn3u67oG5bJ3U4E06Zvi/1W1Jqqbmc+yuD88iccaCEyRoE7yO
2DCPQYJQKl/e7AdVX9Ba2DpKVh2Fjp7/9CyyAnx67NI79mrVZ5lrCMqZDCXSkih4
TedRrwS37epvjZPrYEaCeAuNuIDh//HVNIe8IcdGk0kGzAOPK5p77Wo/dKOOfxoC
ZuBEV0v8ISX3VQs3d/q+OYrK3satnEUlhg1rotp4tIcUbqn3TP/NOSZryVCidcqw
GhGFba7/Km8f4a46VkfVwvjl1W+xWuNOEa8ZdRVFuAqjXaBbnKE+SI9tp6StGXhl
7rI5msO4JCgz2e27dAvEoLK83I1/DnNUCsNdQKcszAF+IjbhHPqFcP0VFnssW0ol
xlcm/sUocCDiyghxjnxyYOseLv6dy0n8ZnpNR0ZItVHJQLiBDtN76T6UFaYdC1K1
OiwIPRgYtdGK/hDyl/8iu1YR2o9hsgrm9Dp5hbCD/e7G40pPKaA56PZ3yFBs/R1F
hXhcPClUb5Ansh2XKQ+JWqatZTyadHKQoCXKdo/8h8ax6oH1ef3XK/Y/98EIZCyP
KnPxkAAgB0JN4rjIzrkztJ+uf1DArD34oq4WPw2NDtRaJf+C5pSnhMVuHxMsssa0
Yxclq2wXtZPpwTKLSR3eyB3ikkzoAGjz00QdOUeJy7D6HSj851pNs+XERDQ9RGbo
dvmo935kY0uHxQSp0YipOQsco8SfkRDdIKNtQVtvgl3C/PsoLoYW1PwfFg1p/HdO
e3qcvrgwPgj4zZE8B/rt8qFpJn309ECay79a3CBuShQfYeCJONVxEzYKYxcweW7K
ztV/XBGPbgUwKH9IIDN6cU4CSzEx/c61sRg2Bh3otKf5FP/1zdsgF1z3QVRTWxp5
dCjx7Hl5yIGKOQQVIgKvoIFjF9t2vphN962zSFpyOtghMaIddFoMMokmwCHOuBfG
QIb6JJampQgX7jzDoP3JB2/gd+ZxUvqEgydAY3W3vJ8EB1/k4CYxy7mYxofBG3bM
vl/6Zc5HFO6qYuxyy7Di6Foj2okgNpH8lFDR3k6tr5rLS2vdMvuEcxqYSyV+GGy7
uiw5pcDgyE+Y8ALj8YSTJa+B3HuAUk2oQQe1w1egmoyCDwndW8oN1vqEdDj3aC0G
S2dnZDmPCqMXOv9NbXqrsxaQ7uqKU7PZcEa9D7wML5brQiHn8D6BHziY6IoitrKw
/V92fehWtiyKVUgMYkTxi2Ls3NsU2bOSwdKRkDi1swxs+Z7XPEb52oh2XrEa8HC5
Kf4zIPfwQuxmuii++PqLIAQkdThrGtk/lNQ9f4HEeAeDKThLxv80saJwVIAmf143
6VtO++UbWS3B75jX5I1fsvLh6p7LCEWkkOvZAXShd+LIZBXx+GGEXDofA1QUIrdZ
N6+ROK8IMfsmLZnZ4izAtkv1OOv/sTNm/bc02FvT4rFdxNrkw+aKulbtsRwgm9nh
GwsJP+hagEFkVK9yMeReLt/VlcxUdboI/ckw4fWmACNBpBwj/rznwqspG9jUpab6
mEy77K1qfRBWWZoKShWJT/ya9gcacRzDePHvppmWHxO+mTfYxNebEhiv3yqRFqbG
/9+kyI+6dcHqlarrHXmWqc3GiIPUgf1QS4MXmH0FdHXByI6vfibKpDP3qydTHjlv
fUUfiBW09xW1XcwuzORaoIKGAvUsk9i8ZbgZ0WWoq/5XMFfKnF4i/OXmfqRVwUNu
9jzJsIT6oH1FK14mCW35MUqoVSSN74XYlKgAcKxcKk2EytZbWzzdfM8vPIGD59lG
J5BSdUiuy6LDgpFyq60w3wfpWcMA1IXbrn7xATX8cHT06wQuPkGMN6+nWDZyd9NB
9JJmBJBPTRfubcywcK9PE7kOoasrdhTl4rsA3Se+XkDLD2i9c9B7IeXuoB77Y6yy
cJIBqmugu4THORz7HjMAUOmIF1nlvOsR5CaSXB+5rr9ku3Czb5WY6x6yh02hVqNx
vp6FKhdGbYB17nOGeq/W98oZwHoWJLnISHKMpe3iGTs/yIP/N+cWGYNUlME31lUc
DLkW30oBtKvrxeWG4geEJgqV9PGuG6nMRiBlBdHWJ4ldfAJPTN5x45he+UybM/gV
V/jZnDAC9wRK4Kz6CYnUf651R2NDT+oeiWM9wMePM6xpKjdJpIvXqy1bT1mimj1n
f4BUuIONpbRd2Yvr75hnwkEhbFy6jVkBOmtPJuSzWuESSMQ02WjrEEG+F99fS3/d
FTGtAl8GxzGuvgD6K19LVTocI8brk5K7pkagkpj8QUerY7EiziI0sAMFxut7hmbZ
b7Crt+cLxhs+sIHEFh5i5/U/4etLUu/i73TTY1SWpfEBePT30x6GBw/5V5szVxuA
ldrxeftLuGMpGP24/8kQrV9DR2qIxdIuNrppwiad7SGlaO1+mKJkPNN5fMS3rwTF
02CDR4m7lrPHrC6LHBCd/h+H3T7ILaf7Y5lr+iytO6u6aZkSeMfgYqw11OtxzUrZ
aQnnVnTHQrJv3KXm+1aasVb9YNj5eGogqgV0mIpB7xXn1npwb1wUc9+9ogvdOvkC
xVmI0Z8RfVmtSyFaBGpOCU3Q9jmxNZbRW8iE73O1tUEUa0X0KG5J2fHZS/3UTlmW
EOS6/fcY9hAygQOkfhJ8BJKw+uSvfPR7D8UkMoXKggtPaGb8GyuqzdqorcADXz0v
GgmUOQKa6L/WIWjB2BL06BQg2sFXH7wpHNcZxDxVF+KFcePXUSnQhTLY4ZCLgV2I
UT5LGwgN1fNGTk/X5sdQ+nDzeqwnOJMnEF65p+3PohRvQFnzylFXiOase4MCI7G1
UX5/T1IIprH3OGJPeRQNZZ46jadGAE2L62gwgaBlGO6P4JU3izFXixgV5vVXZdlg
Mi/feKfuxsW2whKY5K85EMTbzAj8ykKuL72WLGaIOELHd8dT0s2kLQb/IlDiDGfB
W1D3lN3ADt7ghRg6Zt7E1QVsWOqkewZPhPShaLQBqehtPmCab5haeseZ0uI9dWYH
HJ/4L6Hxp59QBmvB9nbhb3aEsUFHuu0lov9z0kskL5aW+EvXcdQcZYRoqyz8H6KE
U585yjer6442MnrS2n39YThQ75quwSisGI/i0PW9bu3zjK2GMiN3bg8Qr0bz+zNn
KcWY+zGho5XrMn+1Ft0bdHYlFROs4qzr13WC4wIxpa7alP0s6zTYWtmxvUjrJX68
QrNnJC2WRgi7vNhvbghiz5JgfqceY1dgfEFU1HP0BslYBWyMXF+R4wvS+8dsedn+
C5AvS1KL60eyK8hyAC6WhcM8mqEo1+Z5cyuFfjHghBnTjgd6exX4tfPIVDM4DAFg
0tD+hXDMCN2gRRy55A6Pvrh8tqun+MF391tuzqaOBJNUWs8lEqYaWN9RjO0HIFGH
dqWbwF4AchbBW911jupD80zZCKxBdgh+U1ubrPifMTMaU0LacelmStuI/iqQrN4e
LZEpuSgw8iw71Yg4spkSytqOZS6He6QPmucJKUVuvwhXXA0Wp2Oz5J/C+PlWyZcW
FQXPkjHODnIELlq11J6auoRobnXSbWRy55jBi3kUMOw+Oz34/oxAKQvp6LuxSbrx
kI/+Uts3V7n2NFuXXX9vnPZy0AqVGaH8m5aOG+ZCBOYktd0FKFy1l1f6QJu5iMc8
fylvEcbPtmBzj2fehQirFqy9HZBvU5Anno7Md3o7zCYLEAlzgI6sjU5vpBGr4wG0
ElWaaFhDRnhzzT3ameN27wTbUyYOlMBbbeVZk9DfkZwXzPsNUbKjNOSJ0WlBD9cU
KePZVWlPvxTiHkZSbAojDma8aQXC77QwXZGXBiYOJ4pFz2RoypC8PGE4z1pT5Yxc
Hf6S24woArJhCLtm8cpEXc/ZBLLpdv9cMa/Masz6bnmYK2oMJOT6SIY9HXB5e4Zu
dslRB/k7zyBRgQGKFLRUjjV+VsEyJHzO8Wl7Xs89kYIqZ+O08kpn4KpyWNFGD6El
MhmRxIUDAnUp/cqKGr8/HW5XzqAB2xPJbmdf5RxF4AzcMJNGMVhpjaNXRF1N3rbB
+XfurSK7/Tc8vvH3Ggcl9GONmGisrIVL7wcIZweKZNwgdzIw+IYpeGlCFH08wgW4
FrvS9/IoarqPgxowjKv/heEWV9icMH/7MuaWJkh6nDZJiN9EsV8Va9qGmw/DgwhP
UOOulKjERwV6KC8Wz0bzhun6Yv/auYaG9t8DN4PSijMcFJEso9+AZDWUe5ZlZ5TM
uWKq7UsqciddqH5YzeML4R6M03uLOaF3mrPKzIpG4h+AjwXAorLM1A6lj7RCEaaL
c+IWF1NVm58Hs9Y7ef+mOv1vHfg9ijoB0SkS+8VgoIxDGX5EvUSVkggzht4+rmb+
mNF74HK9WbUe2kA3+zhHwKWmejHE4OoY+m9SCMzfxpkwalb4pX1o4UlQftNwL/JI
2zqyW8deuO1TgcaEiFVEKw3MNCTf3Q1OdcNMgoK4WQapzCt4FqmsAdxPg7juAcdO
Sm3RHODN1N4acI1Pb3CfoJeZxCYJ5ik0qtiPNdxfV2q7kA9uUEqlNgeKSIEjDwAm
YAVS7Zde6o2VmCC1XQL49Icb+XGCVmEJYcsgP6UvK9+AhRcliLca5Ar5TtPMSU2d
/pEbSdzXTLC6LGx9nwQY3RN9bz3sDkgHdnKSwvmL/YkdBfODYfYld5VlnwVidOcR
vjUhp+bfdu2fSreyNYRg63p06Hr5d7ebK5kdJy1fXpnWQm+1sa59GOFcizVy7K4E
dPdIFoACLm9fPt8/J6ffewCDqJmb/cxowK8bOFMf2PIxi6ux1oxgjY2piSQkD2/9
qWWJhL6dYcBFN/VfUdifaPA3+F9lKZJ+fbXd8na6SXclEQwdgGv8Bzp+tuyxDAPC
GLAMbC33IkiGBtZEUL1c3DP+IbG0Wh+I28S/ws57FAj+P/vHgq99oRv6dPSL0vID
QhjnepJQbdg44+7cwnoQL6kyrU1NGe/ir10UpJRVG8/kaA+xX5T9BO4fD0PExUat
Ak1Os/E4aD7NvIvaHvUSj6lCNFPxacUAU5AVCHCCOUWTiZEtyT3oQX7aQ++5J1XT
u8LIPZpvjgHSbiJOiRDLI9b/qwZhOG2sNWOWsXceuY0YFUQEvQPE8/hhfGUL7V8I
Vv93tcZqvm9XvLlES3rH6sqlN+vDp7GJFZc9FWI2hiFukE0T2BqDIpYnrm18MXrw
Q+wyIqLvXs1HpuWCz52tgjm8BH/2mEX6t5gKkKQ4rF1yAqnOl1JpXEVPNGVmQNzO
X+isHluvzs8rfA8Y+EzWC5gPJJRItYuE0szbhp8IZQ4uIxXRTbhuOUnxDLfNP8K1
l8rVIP/gy1HICJJrNEXjoKLv4oq9hAqwCu6LPLuHs6gnzu1kPSMQRVblNTQTjRZP
xZWLxd0P3ng93NVlGqeTDEYkFnFDDLUEuUFMDLevq4zZMrDBe7WfEE8OKwUlfF/k
rSKPym4eEoWwLakMpmZHXfNFHc+DONCByOTK0vNlt5NfTPRxrsYtXceRD2HdwENr
zuKeOcBpMk0qe2FEb7qgoVnaWvrx5MoMcO2ZvC6ir9nd0tAZs0sybBPorpIKRdIC
JecI3UODLsNSZb8KNeM5usrofHeTIZAAO4kREJIIGp6jwr59+/Y/hf94AbnFPIt0
oIrcGgG9hwkxVBaISzsMI+f9Y5kHonLyBTN32BBJT3toK9MqRdqbUTFD2niYF8Gq
zmRCFobaYemX5jxjdLNEdJI+teEwh7vtU89dsv76MSqjQrvp5eWqzrUZMHvImmB3
uWd8TaQXGtkyCpYjgkk9wKFA9gzXBhPuyPNnNLJQXAmaEJ7Gnh+xytY7nfrtnbgs
BIF4g++aRsIw8USh/eO4NVySCIrHxJTLS0R0HGo1seBuPb0CBJoWHCXRyd6lign5
rKtcCz0Rp6EuqhvA4w7xSGl3SwmBwxKsGzVQBBjUxYNwPzwJkNzObvQ2aWX60IxC
3p8yoiHmJ6Hye+YpbQasqPvYSowzm3llbfcO9IS9vzscIKiuJ/qXukI4BoKylkMu
6z8HgtefPkTk3Pvp41Qq9LKkdestMgwgSL7XUAjCWP/54pCVMhg3jYqyhbhoqNf4
dvZtRszSySnfSyOcfOwPkU8vCPDuqhmeMGqFt6ILic+Xqdb0Z/i0vlRd7G9fbXZ9
aFNzrvidjX8m8p46buXAoLf0V6eai7QDXS+wOiQ9T/0/RP98+wyNba81C5bj1326
QCy8y4v3W07wOcLZpS/aZQz3q1i79a8PS20jDFVsSqNv9kHb1zYGyiC6NNU0PyR7
0sM+/nDSMua4jt3JqxOwKCmXznD3H3fusKYQq+dTOG8RjD9IvS3fmObP1uvYEtVD
D1sn2mmq6ZLGT9IGRclOQ2jfoSfMiG88lu2NGwgTK5YSMskGbT30pu/Or/69ldJ7
HguRtxsTFz27hlEQspKfTHllSFw3wcPL88GwF0MGXCAQbJ8V3UTEXttSQlkz5+eD
VPMXn2Jr4DiuLvXw5p7OzUNiUqGmQvDQAabDaVkq4+veoMBExchwunGyUS8DKpr4
me6OdZvKHckc8TfTF2yOu7qcUK3qCulcqEzeVO1NQtCS/eIBFuE9JnAtNUeV7tFF
6uyw53b70dUPWKpfdjd/U498iHU4hE0Ibi88lxsZ+0lUTfuuXYgn/l0xc69M0sub
hPPGe/0IwMyedgqGawZXKRSWHcy8dvFsFzZunlOusDRYyeXFzlfqLPUrYRDLuZ76
R3cSMKQar0GdXzHLzGIab12+mDq95ICChHa3iN/72moniUcZT/QzdWq1lnjKrtkJ
Z0yoZ4hQMJZYZCdEFvXN+Nc7XpazlG4puHlxdVB8k8Qk0perZfJZ4KXk/K4mCG4a
LXuREl1GmtQ5+gJkXScK18ef3eZemUgLdhgeRnxhhKlkPZ4zQWyYyy1mp+AzOTWZ
Kp0CSWavPspHH7TQWTb82Yttp5Pnm3YccmoJXEisb15SKJvevgadQXcclIiBtMKH
ZocKfnocx1PyYom0NOv57eItLGt+KFNdZEqLEC4T13na5gr+ddVEa4n9uQJfczLM
KKRMG0NQ7uXKTw+mGQ9AxcU68+tvNt3FQm8uehnLgJmnec/zPwon6lbveLloxOLI
OGFhoiQ9prl4G440wCbpybLylZx8YBPR2XJ1WxxxqWmAAhgrkRuM7a8jdWlKqpdI
Z38FBYYP48ylZVOv2OnzphKvaVN8msTCsoVe6jhzJPg5RmuF2zNHKKujxDTB94R6
joXJ1V/zlfoeyWCgQpL3KeX/yEugeItgHCokRf1hdOaVyGooulubty7chUG/8Pqw
NsdXyt8ofmt7oo/EOJqGmddtpe03V7p3vgtfNwf0L1RPaKyc5FdEQNQMmgF1UNjs
SxDGZpGGK/80KX5RQI1JgJt2YBhFNcFLvOJ809ioh10oiKUkU7yL0eNQO6+tk3Hq
QFPTiWFBe5/Ud1CF72BWYkRFEt0cZ9h1MPndPVhD1daXn67AZpMNKTUyRbYjPpT0
ggscgIaKiUy1rDHB9ZPNSdo/zsfMeD0aXATpyiEXwIcO9wCAWDSCgI9PKlb/9055
yIXlcPzjOsFYWevk485rpAO+K4CbD+9/lsaKOw1NZXVCteN+lVUKWlvDLeFrSeA9
g76Oe770RO5yVxb25GpDMXI6KQzomq7eE4xuQ3ZMC31E1Vopi65dbiUm1mJJBob+
AwNg7PPQnpYr5CLWV0nv5yx+xF4f5W08IE9QvGmUX3VCmfa1omeK60HRVRrkdTQ9
gUzxWf9PKF1l/z/EeQ8enGFy9ZNLWrUVWn8tC+XRsKd5CoD3YeAXSbx2FA1ib4ko
QOZwdnn1OteXZ6k51yzaNtIOpFEPNCZs7OIvbFr4ImwwHM9luoz/DdRrgTsms1hZ
Lf0sWEEZdaqimws2r96N/Tgu4KMBlBfw0BIxoBcLJ6Z67Su96okSYaCBm43yi5yw
jOKutIvlm43jXd+rsj/Kq9dEUfBuwFpJU/+7AYFiLFM5ntFOpS3JMKb3O3OVPB74
1KVrrVwigxOrxDea05blzG4FbdNmRju3vrAVECPmxZ48XcGNCa/Qn748HxDJXjfE
LbB0y4wiTSKR8O4kvMZPika7jD7LnBupl3RiGaSqvXCCNXp8XLrBoclH6Wq1meIk
DNb7Sf7MGwMYwSUgxrn+7ofgKrrJ5M5HiygsHFSAxlbWlMY5NPFthOllKCDdF0Dh
6idMHPkW8z6s/n7dh0X+sd7K7gqaROwyaKuzRlrOVxl1I2/F29++5N7Lj6BFID+4
fcdysA3lbjUh7JO5XKtPtOAK9MF+IHuobiF5RsEfKaMIckDKRehGfJQF9aGkTIq4
ctxoc/MWTckdKme2kFtTbb9GVPreA9teI7h26PrDJ2epIYB7Aq5QaCk/v0+t5NMb
zICa9dOvlbSAMqz+/mDVen6H+5AFQ/dF1KJBO4kuSfuM4i+tXaxeNwDUmwUZmc9d
RRg353Fx/MsPuorsVMJZOehYofylBd+YHU+r03Tma3TqW9loH4ZwQTtBAsXxi+zI
tZaZ5zt2lpBWa6ugRk3zd7GBlTv4I9m1Ufct3N+VbSwFeleUHDTh4cA1XFBooUxl
ARgXlPuB74ecd6Bgzwp2omLulKbHQiY3b+jYAiiFExP0OVdWSzfZyMLEKHTfXoh3
jSuIxjuLZz4gd8t4hqZ/J8lIRNC8aY6o2UwW3/6/vSo8wrEVz2e/SpanrllxCyWy
rfsDGCELg+Ql0/RfN222h1CT/vV50221jbX/DJrcX1R3raod4tGfvhHAzELO3RTC
P9vf/+zZ7CDrLjXrRc8BqtEIVnc+FpDhwvvZRxBo0+/hxI/UnXpj276nzNxZCLU2
eFvVVvjaB7izokJNpsfTMZxh7xYWCso7wXNq3eukXjAbr/Spl6640THGWHAsgTF6
8/bMfcIQeh5fARJvIhg7veIqF9uBApNR+eTAyNlk9gHIdaWNvdNrCsSOw1C9rT8G
dLPWQFSoPLIp0i4+VvP7bDhyv9TA6B7l0MrBG86sDxQAjimsATF+WRi/CovCEbRE
JLi422tqCi6prNf0fsXDRMCCbFxnra7V4X1z7qTCRjDUk/ZM0fBzeQBazWFq4S8T
JkZtHOzCiYamnK35DP8UCCm0YrTRZdaiTzv9yYKvO3L1cIOBwzAmAn3e3acDSdiv
Lyj2CGJp/RRZnof8nJxkJcvf0WFlZIwQLyP65Aad8tsD9N7YdgBmJ8qKRFqLyrNq
tY284czwhK6CClAou86uv+wUmvozYXzhwJMRbmjmBL+yuSTcsAq2/xMc9/qsHM/u
hMF77uBfvoe5oyxwnfhxCWS+OE7tIrXJ23La97u9obSyWxXBUU+EM38heH858X/O
DyeIntnGhiITljBLZZdznj9NJ58aXOhhwwCcSEcYVYHgf2oLd1IJETZfVerXNV/m
vZ6VoTUr/CJPe2pPCxBzF7dVzNPj42iPqwm/1ZCjN+QiZhSi3lezX8Fa3YMlUoL4
SXVBdyfBAAmYSwMvqjK4QixGDU8K0TKQfLQBjVvEtya6zDN6VO/QY6nD3Ix6XYbk
wjB4VAQX7Ob1La9xjcLw30kjbLw/Y3t+lsGwtZ/+yIUi/eXoObQZSm4hD/fnnVzp
y5wEwugaABifPYlX9icAJEtsOuDjkEMo8/ThBpn4HX/u/u+7imPRJEuSmhfLH0zD
NfCi0ZdTQy/uMT/ToWbZkPYopv/bP+hBOzRzvVLVljL1z6kcwlAFXyJ46DbAD/Rf
NaCKfQl9KHaGbcoliyzvRpRJZHcnS9ut5rLXys8Txd1Z7eEoT3Cf3sUgu88Dax2Y
nfHgiiSEiiL6hDXbyRxp8HQrX1UBq6X885TYMtGJGCQAifgp+Mem4jIPmew5//Lc
50G3ArF3LSFxPxet+DEKkSDe3NaMzuamlTfuNIJ2cPzjCB8qGj1fQK+0TxOFdeP0
GP6FHlBmk7Fd1Wzjvfb1RwU/CYoBZ1sac7AsaSwLsPSdmMqWBacYP2h5BuKLWrL3
ewMzhPJoSS2klbGYv6tixUeXDBBK5tdctbLbY1IS9txSXlLSDnrM04Fg5YSZ7MiU
7eMbwty/5HfCc0nOHlyp1B2VpgulrcU7t+4NYGlZlWJ8HJrilyF4ReV8AKHlqoDS
0Nzpml3w70CaE7LAON6a0dBOwjjhUsUxmm/K7g3kLmQRhnF/qa9Ovvsw51tNEDwI
mGdydfGU/Pz2ooor2V3QW1yOfn48sCzYARaDF+MzaFXPjSqq3QVEBqjULwP3yHjJ
PQdOdqFjVgg9qhPL/m1AMBbQRKLOAmqYZSwFEiBNuisjt0bbgQSHRlUphM0QfZ7Z
4Q0aQmquXtURpx/75TQA8UVCqYcfyDZ3leP6kire6DqNYYLgI+SYVwgnusHeFkJU
oXdgjgLJ1b145kf3eJn5wkrkHqu9Us8aTej+1GTMQwl1FvzWIEBzAt4RGnPWLs4h
4kMdg6PO0juuDFLQN2jM2wLPj5d/kynxW1ujDxgPCoWr6XEGXel1P5PLTnJK1kSx
meETCRrEFbhUDKB1qqE1CIRlGmGNqWUsQpzet/qwlU2IiVPA9gzy/9z3/fLtry3d
B1GtLK3KQ+98m+gCAH8Gjdh5vyPiwI/0ZoZL50nfI8VVwzAIN/OiVWlCDiFi41BU
devisLWsuEkhQbFU47EItAxKfuMvG2Qk4UfemD/1KTCqdmQChkqx3Ox+ezmQIadG
pulSSqQu0IRwK0DT2IBvaMnhbOGqh1VAcPO/JCqkn3RLpbm3zF0j6I8Wx/9rZZXM
0d2CKgEuPC1G+u+hJKcGhbnNzLjnQCsSlb16gcI8r7ZmWJc2KQxT6Grep5wWIfg9
HgFAk4PxoWMo9lTMLNlh69roI7CMITkDIOmYSpE9sT0UQZvTLbNj2yF15a2/klFU
DTczJxB750WGlp7X7sNxw8lryEW9/JonLgI6MQOoIgA9vKggxHTpw+upEWsIU6hn
BofspoMvDvGB+jIwnRCYIHXTftlrFcTtXfrPYJ3picDMGJn9Stkff5tXCbhBHRz2
wUApCZPA/0RlqdvHHaJIBVGQHk195sVmxHvziD1rnGd59xP0LfqD6uJ0RoGkB5I8
KxQrtDb09G29ExKpmSLsAg7N4eCRKX74VIz23+PSxS+IGbyyqNfa1NXieppSVydw
DUykwOwSnmbR6oACkjI+ZFOLaH/+Kfrqba5oFvAagngxgvRLg2aFnYuCbxMaBbgb
IGYIFxt4GR5/Bav2bONrH6IZ9DopC+lI0+le5ndp/O8qGXHd9AtrHazJ7q+KGnA5
epoTpWbH6iKR8P1oxW6e6T4Vxws3BPYK0a1i44mRbgr9IlhWXoZLGacal7ogPb+w
aq3edwjpLd0SxgSZwe6ibtQt60onh/v57TPkin16dOA/fSRFrQ7XPFmqcwTlbzkn
qFAjzHamhAFWeipq7uCSXvJ0HegDzjkIiNIC41Luj+9O3laY3OIAiSjtZciacwBv
eRFPOEE+2dlzi9A647R9r27zmQJHh2k898/GhcmqGfekjkQcL5PWuxHlOd6ko1oE
PojJYzSKihYwz6tmxWafZR5YzszU8lCUbP467Q+7hiK6V16WLKPL4uBRw25jXd2J
qnfT1b8exy1QKkw3SUnHSSlpiESYsqkeec3/aJz236Vv+VNKxsdVFcb/1nu9wCiE
1svtzsbVQhhgT5FY1IE+WdKOIs0Hs7h4q0PurvYiuKiXjEmizt/37fgVjiHJ/+ot
nIRSoDT1IdNBi0vTVQRyPEZuCKKBbs2IrZcrhitbSrCnfFMjBabHu7Y1BkorB4Uy
LIoE6IGz1gY25dZLjkpNuVomzUHJq/8n+Y1Pp29uu90b2O/wGn9jqigYC6tnTo4K
bhUf+8tHgAcwcTJJIIpHU6Xnxb8zZaXCxfBjJ2bDd6SjL9h/tRbOt9RULskxw6qf
2C3oYU1JUmGNt9F38+ArXF6uIfMgjli/S1y2+tzSOzB3v4HMxF9aAtsXGFpBj6zL
r1yhXfwcO5PPzLyyygJ9/xIYmqG2W67ayxgacHgq5usnBLBkS6VzYnDTAwYK9cQy
tFnCDTWhjVTGZmjXPiUF2MEYTM5v4kQPBFfK6Nla8YsK94W7TObjuC31qlR8kljU
8PBfTz47HPVgd+IosNJ9yCsR6zovzsU+lZUqsw+B6kqU68DyIXkkNH4MaVQL9R0a
qrkV9CcDcgT3otzxWyObi7ttXiW9NiroTViIT0nxDOrZ9dIgMC1J1R5Jrq4gqQkT
Nxu60uYhRozAas4BHSn4ykxlzpRy8tz85tt0Iy8YFycxTuXAqRvRdpkXpXpUv5Gt
smoY4mtrWkr2OLg6BmXzucIMNxsgvTTt0q0f9OPn+QnTFnGXwIFhbioN805lYNtl
sQTd+3F49JNyaV5V9CHW4PJwBKHe3szDys4OJ7wph28cUvLRvGipvclugORSnkl9
2/kYdiwDJzLna2K3q/C6CTlhQUTYRhHA7tSjqTsRjBOc1wpDoae7qO1Wo5EUbnqJ
ttRoswx+T3HZNAn6xKjy/qOOQdq8qlRT53ezs4r0IpNPLYQ2CsamC2i2MYwEPuhk
416qfiZoK7vEsaYHJLTDiRZdktopU3p+e7geed4lFNtuDFhQGABOfi7ux9iwR5bs
WHkYbsPnKOMS9r9FAE23oiLXS5chTZURbKcM5pWpV3Kzv0W9ND9RVjLFDf7I0tki
IsKlmX9DCJOhuCk9kI3gW+ys12eIVXa+mwxr8hpiubr6MAZK4dG80tPvf071I9v8
eYCTt9S8ohjdN2Hw2cDE6SMIjbuJP9EG/CnWjZiAQS4RUafcuwuyu0A3ZZtAJJxX
coRZjiSWk5CeomreH2CciDQFzjWIJ+N/aoUdskiGMurAcQDakD09Di5U80pGTQKw
iGZQQZ7b8tqbmWQFSpFTQjOVp5jgoVDQECkyWLmtvVK8riSgU93WsiyFtcZxnxAE
E7VSJtGYQibPU0yQriP644L2Y1cm09fDvcIcuJccRyrGBcyMKtfr9gIcv566hn/l
wgv8DX+p/bI3doQSV01pcDmDTnj5FLy7ix/jXLegqOdQrJKdCPRdx3l+pL+wiqLN
+wA1gFWrHJQIxrW7ObX0c5sH7csk9lSrmmKe1J6lqP1anYndA+xXw132T60E1vs4
f9ndn2FarvvEHTHxagDsbYdbtx0qZUcO5xdENWg8q6P55++e8ZxK4r8TkREKeCtN
BpQKLHhSH8EHYk5ZmandpZE9a4+rTIQvZCwtUg2auad9hiqkId8KVgFo+kHye5zX
rfxHM/VjrH+vZlIFf/lxyXq+H4JTsY62ruhlibJdlEPxBRw7NYEKGK8m0gqMxpRk
kfcG3+0wtA7Sbaw++h8wcNaRYzBsQP1f4wRl8OnKp+VnXZLwP4anxLxetz31P+Y3
YyhM8lCzNAt9PHlJBHffsvhEJeuSO0np3i7LJrf5YjncCPpQTuVb6fG4wQM6dSJi
fuMfSmIvg4b/TlJnp3sivFgGgakAFZhY2qdqAjU2Ov+80Pi/hXHDm237L3INCzta
6UJaL+VpxVYs6f0zZNej9L6+XtMJjmBXZMGTwQ+0hnp0tWdadHY3t5wL2LcIkNm5
Bx4Z5f8j9oM6VaZlPDvNQHXwZEDgcyoKCmr6U3Wfcp2/8Zc59irbTRtuZscbC5/w
EEwY/koQkPjhviXBkeqlC/DUEJjkMZhYbsmgrO6BhSO03qKbc0ZO+pujFyu0I/80
LFD7ET4TEhNscjd6+8Xg5KojhhOzKgz0rBVROmQngseimCVs2+VJqwX+YweFGWPf
rbPqqbf9ombQChnkMeSmMVmfJOe6dhQzffu5LnA2tPrSB8NmHHP2YtDwfaojVS93
+BUVuhUB7KNkNOhP9K5nvkyqnOus7+S64k1uKE66bhEqj4LMXXewPJmWfuK9CK2S
UowR71VBEy3eps6aFL1QdWPMNw9cdp5tGcCOK+qbkPbSJMN0JIaTGNOz2CwJEvqa
TqWS2BFzk2GiZdAQtYVrQSTZMeYkt/Dq/TS0+Yw4O5TMQ6vEPxXOEukaMhV5MS7X
0ksolNDEvXIWKpbCVE8+x9PQnQrU2XY/gZ6rNZRTf8VIX6eoNoHm9pUvSpBNsdSC
56P+mN9siqA89LDhWImJCn6OUb6lxRvJJKhuoGQojdvMdtzRBqtQaPuzZ5KYOcmu
nAm5Opz68rtdIdyY3GIdahC6trcHz5n28gptR5FaIq6EIKfOzP2A7+II5CgRiqGt
m0WS4sXQ2NHTHO61pGf+EClSvLMg7naFwbabpUHp3sx0gYqWPs/Hd02HCjCvaTiw
jx6n6p++fiLcN0PwzDI2/avwb4RKXSmXk28JdLWcF3PKDVwuJZ3n69v25rfzn0pC
mBS9ZNFMuJypZznCf1f4pDHLawUdpsyI+3YKPliL7wT0ycK1ei/uA8g0qsBXHz0l
NuJwuLxqCZy88F5ywo3+P1TsBkGVps+YZPdqdyrXxW+KjK9+yTRn7XLBLRgoL/x5
04SSNnJ2M1Wm3uAJjKDbbLgQqwFfzQ1SPwHLdQKnn0VgE3LjwVLCq11Sa77RMzLr
XwoqZl1ck4tJbXHY/JLELHOvK5RdrXPbKdnrncEA8cKwWe5AJOGW9pfo7RaZ3siC
/cSm3iMC7w2lozYEycnI/pFDWNqOle1qO4reWpaVUczRH0HKVZ+AE1skTK6UopO3
a5p+jewf5CsrYYfTlrZz0gU/HqVfq77n9h8T1SFC2qYUrjX74kJ6PxXT+F1155Ze
iCb/t8yLmkQfsMt55KdW521WLnY7VpBhAsEHWBP2wF0AfwUYGhVIbvT6BcgA89lS
7VGaC51+uIfDtvtm+kEh1j3CUtx11/22lt+yQP+G97yUjKkpSEcJiLND2XBdTdrH
yDYbkdydoY6i+a0nIHC5aqNPSfI2rAMq55KvzZYXGox4GAb6zV3AflSCfT4gn9AY
9f8U7sRhWEURYkCfVd4pTIUWM+zg1nxLsp5K6BlYAOLU1OJDgBpeU5UiRylfsD0T
HU+0EmBXWWIeq81jSecgmWQwQh0WPk0+Kpv7b55oXFAT6ux0xowKwYFYtYKwkUdY
T0kV0SMxCDDncyxc3REAnVxJN+YlfyMRgQ0pPCUGdqj2vnUw6/qsgeO4Wp7dBhUU
8dT9oFxXWErILsrNrb2cZoCFQw5M3Os/AH3kQpxGFNpQS/KtZEZ5It3jMTiLKB3P
KKQi2wnYp+W1R9D7bDEx5sJ+0C7Sf05WDnkOoVIOfpjAVNmPeuA7EMh9ppQLvdZO
AUuPcA+FiW8xyCRtx7PHwUuvhW+zh6dwlDQ1M7lkd/rrCRmxa5DNcuFGQktCFreD
MWOowwzd+LW0zhWQYzPivCyWCpJatMUNQSG5WwWB3Pav7ipV6249quFKjO3o6k2Z
/xgfUDK8u8KMIvcg6t5wcwht2LhapR3GjqmWMVaVPTSjULwZPrnGTqZjA2dJVL4y
G6XwkOjDydonCNYKBOBLUpm4TDvPdzmZhGq4q1rHwSOhr5LWL37ipVM3DRtVXC3x
46A9/w6JLHAnrPHEIKA+ceKirOVjiaJHGbZGDJYmXQQAiCQHgHrlXSjQIIQ5wWaA
VR8hsHPXDG3Qm//F7mF+2/09qKmkCHSBVa2A+WnX1aouWYuG5k98o+YugE+x59ty
KTl2MruvC5K2zS3J8UL2PjRJp5AVWxvtyNDbczJTy24DukwhFVwIwUBp+4uddydY
QA9Vt5dbznyAmsrLb6+fCUZ6jPMYACixAzKZqdAOOGNQJwLlhHwkK3oPjIWdxhhD
eEMVTe+rZCTZYCvKTkQdwTaDanStGaGoxn9AN/XZf6fqWQMDYtzy+PKasXJ19Tzl
WYHcwTsRVsErEDLlUVINILrodPFlNQ5OQvC9V/OQ9stDkN3jQ1qMaXGsKPXOZkA0
lP+9aeM550j51ZuVA7S2tZGVGypMgsCqeEiXkS0ieXxNFlQJTTWW2WNX/SqAxXNI
OI+vKWioFuPuhkjsVsmHey38OX91IlXX0Iogc7HgQTZ7gNcu47Th1Geg1/+MM6fm
59JVpz7VyPB5q0EKwu/lHxFVFjlBi+0lcw4Q5j6XNlN7f2dvl4wET4STSChJLVOs
WkMGjxyyz86gmIfyZqM3oPlG8hGgmXhN+U9zRiUWKsmHtlyew6Y58BSS62kf8ADJ
JO3sKKdC2xQ+5rT83j1Vbwa/0fGzze4wA2gz545vemElEmrb6B/Q/pxkF8dc1CvH
CmQdbJf0he59raPgxkujIKt2+HAvx2zQkpDUnDEEZ4j5lr+2TxdXvOKd5Jm4D/7j
LvPZ2lX//B6WBExe0FU7xpAAhu/AK6okTkR/xmcpCL3MOqTNFVeAW0IxFtUufpx/
PdyZ61I96Loc/AbA7qs33zVFPp66X9WgSiaMRDlAdbpXershRT1kPqBN39L3dwky
A+tZsNQKoRGqkNv29U9KdUY2c0jWftEhOOHEKc1Ud/88KiHWr7Mcg4TCAj41CKEY
oD02y2TgiyoXBW1Teaha2WUjcY+Ol8zKDv5tLzEBrRDPcV6/wmhjg4yBb/5Ppgd0
sOcUAN9eSLKEzZ4NlumyLOVZ+XY9iiEdbn6/HDj3/aS3InEH/gzJOIVUOwjCosfw
H4uXdcXnk/2rbJYBu+IwMNX1RgdiktdGE82OsJf3zqbdxiOBr8toSfJK51mCAvIK
hgAJGy6u4cvTy0I5535x16Duh9tFJF7ZvMxUOTecflTv4Zd1PDOgr9hsRma9uibS
p3EJ0W5Ywv2kw5Er5vi+nKH3s243deKjOwJeeX9D6Z5iQNOcwk0XFgTg11AhTcdE
5zIJMTwaIqwgbD7CsF4ONcgyKe5JhBf55/VJGde4vAIoOm4OJQsoc0rRJdh0bEFK
LSofW32ayNM2TudRg3IPG4XgE5+BoSkccAC/xrrirV6zvLVaYAHUdEDCV4P2aEWi
vXXSrPyFLxImxSycqsiGGWX4GdkYA8qEidb/pROd+8QeKFDmgGv5V6HQZeCrIWJE
7oi0NtL1L7yF9cCpHjn0Nw4llDARaK8xaefUVjgFT7tKZ+khEIV6IkdtCsicwHIk
vl+6WHEJH9C9oCvPWuI7Fb7J3VdKvqNIUfpGVXGCVGNLs1PjldJyXpcihgjDTi4U
vgchFKR7Uz2+boiIiV0KVr4WtnN2Ztu3XHr2KczOqZ9zrfywDp45NsJ5C8QLCnHp
NOsC6m9xxo/KNIM7zBqYV93WZdK+wgQxqihborcpsE7tjCXSk2EVBoFqwKFfX9aG
eYtC36mkvfZO2coYxXiUWHMowUHS3wWEugluamdoaBa3oprsDqzsktH9PWKNHdHv
BkT+M/9h7gXEK5itnsD4rygdtZ/SRrkhPB9TIQ60ts6QhqWNnD/kmklf6g/1twSZ
N33Os/wLlXQpB3kcUlcgsqBq/ElR1uewMhB0trWvIsq0+oKGZ7OsmQ3nlwTgDUD+
Uxn/BTO+lUd/M5zVa1Ags5ehRcnteCLAWFVvcNEP5i5JrDsblOt4RTuIOldtUdLq
a/Kw5PxjX39+VpzDi3YPY5JOXiXVvrMedSUdyQHW8yZ25RKbQTmmB1nUujUK8H0J
yiGacLvXKViB/RMp1kYcWbhHiTpxbqlK1V5PBWnMcao66FToKtsa7Uvm8IQzrcBx
8G0K4FNSSraZmwTosBIZ8gtha+s7XIQ58bT6MLKHixjBBfZ9+cv1bP//CEaa8YSJ
X1pm3uLWF119UhTHrMvJaz66xysl/NtQkNPjmcpQYKGydQiwS0UduTFlfXQNiXy7
zZBb2lGqr9Nwoo/wpb7a1wdkbKEW6UvvLVamjNmWnlXQ4ojFJH+PhrCq0Ss2XM5P
3jhabR17gNsUZFVJn1g0p/Ef7+V+xhL+Zg5X7B2dnQLpk49gBoQXCUwXpzDp8fQ+
ABvLBF4s/jgPYBTYar1aH/TyoIbiBVJpO0RyWWBsLw7U8OuqqmkqQ2fD3NMEUuk0
bePc0Pbv9ANxLfdCXvBOlof2mXDBaQJAJkZC1FqR6yL6oMADWcKDB2RDA+5DRMN0
6xnrs7GgfY1a4qNqBtVVLrLjjBLm9YZn30ct5S8Knl63bbcPwPAxqdlu3z0h52q5
of0OdR3Xx9BhaabRDWOG9mx1Z2kOCPdC9hqbJkRaC142IpEawZ1TSrpImEwnCI/b
tyCmNT2vSuQznMPAQgAMToq823mW7w9w9p8EjMMWQ4lX6Vg+JphiCG4L6cNQWyW/
6OOyQoskDE+LsWcVL7H4m/dU1p4+nQJugRq6JQxikQ1ecV1g5pqkfi3PbM2io6hB
xQoFYdTmlgLwbT+MrQJXsMBk9RbAZR7nBPBQBWt78+db+0ol3RcJYoTp/g2s9PwI
Qo7a1HhAIbbwBcEga7Z95PajR76kxxLKhTlKtCW41xKig19IbKERUNvnMR6AaLl1
55k6mGgpdxcVMdJpN++TXSeJpUNSAqjvdTVrmDo8bUdVNP90XXS0Et1iUe6ZDPzg
PANhf5WXlvmsVNo/0IVcO5QvjhgP0310ygrDPQapjTuBvac+jL69JzIQyJghZhSE
xNaupfhBiOs/EJZGPrf28mg8TePnWC9gxDdg6EgX84gCX+60QZZ74mvlyOcMH6gV
x576dBPj4noNmK+TbmWUu45sWcBgpxsMIxzhiJVq4evvsxImkgAwPRbiZtg/d8+Q
pkD0SazlJxXr7riSGBi7qXNZPLRnD80TsVbbzaq4Mhjl/y1fFxyN4h7+Z36hon/p
jl7HwlamaFQH9HTnoXQHvYO6DqZU+FMdDt0egLWh3ZnK8UxRx1ZA8kUHXZ1anGSm
x7dJDzL/rrnlpW+qpDoexJhhJNbmdlv+l0jRog/ddmGnGBIuqgj1HrjKBgb4Wx0P
JxX3C4Ih7uLx+wrdU2mY7XmK+047sRyJNkDpc52nEby1jG5UwFF8azueQdJ8Zp49
1nBM2uhoGbDomv+xOA14ZvEWPt3VrdPWLZBJw7xMN33gycEQVK8QozsiUw2HcQug
AVt6SpMi8mFluygZSArVfhP+oPvyEohXueG28Xysy1GTgeQqgTN9eKB70Ooq0NAe
9TwMDe+Im67276nQO0ejMjta8WlYShwUmsW4TUrxAzHGpdK2xCQ3cFTC7KHAxA62
gc6OvyMK6MEi1MZm7+2l0f58ObsyNPl5EmfdeNqUrFQq3eHn18Qhs1T55UcmcXup
NkCMQH5uEjd+DbrRiBuk+JHr8xsEf+LdULo1YKiIG5BPJLhVjARECbdX70PzVeiu
I1HluLrfkScKZmJToekMFqmCYDkBJK3SoIIh+GW17eszmJGIXJUqDFFUeAftfPT6
Hmlqw5Y5FOyULvfUO1ESePCzJy0PYXE3emmdcfzUUSMCb3qsaLHsUd4wq8H8k9z+
KQZnJcBTwh/Qs3LNZ/VtRQFd9tn7htLEfLjXD1GxZsyYG/oyEjO8ddD67yQZRogQ
Fom9KU3v5mACWhq+jH0N3sZDXtotSspGfSnUocCV1kbWW1VZkpKLYivrrIzJbSWM
mgYWZSBLbzaLwYA5h4NHm+EVtaUkrsMajwoTyU3C5NP8SdHkPa/FJu+ahspAI84B
vAqn8w5ikKbqSlLszogn7yb8qdoZDv0OIlnmg6vcvxpJYTwKs2yXlTJQeslRJJet
wQ0VB5i+pkx2P5ypMnAX2WV7BxfIL9FvTSFVZLkSsu1sUMNd3gDI7/3NGKnHmX1f
bS8pgckH9aQgLbUdFLJ+kPOWjrWWRHYVzC2TXINqYF738WnCU6Pj2R08L0ZeKhw8
+bkk3Q09srGTF8DPG3J7ZVi8tqRBIOZJFBYOXzygQcTJUCBSwaVu6hBKFx5T44es
kYc3NsOy7MIyMmDHRLKUf78ii78zp+sn/wD2PMX7ePP78W1IY7dcN9QcuWfTcnT+
GJLsCFhW87PKr0dOk46AAggWZGyZZQnvnRkmgKbDZefz47buJWs8M64d0M2RI9MC
Ld//PC7WfS9t1SMdHJ2vL2Ab8kLUGfQfLEQo4W06JDUftGgMOhxcnzh6nRTk2wtS
DuEBguggEOT3E81nwWsUGb07PXv+YhR8pIpaBwQoeAEYVo6MqwaDDre25CtKKmit
RrHtIW2ynFKqzxXRCudvwP10LgT6IJtORZijh1UB5OYOpSxtUcHafTR0Fnvmhmy2
1mc3Q9mja6a9fBcyRldxBS8fpFvL1znPSYodQwfufnM1VMxuVLAH2hZC8tq8Uut2
2n1piUR29MhTANjXU14qjVa6YkAaaxB+vvlH00ndHx79QSKWOvIKkDZEHMJeLjzU
6N+sHpW+Yrgw25v8jngTEalqzulOi/cFPwFx/lAzlAo7jbqhqNnCdqjkmqn6zvkY
D4lkrH3ysQ+08zP82n4psP8NkEUnAs6EaRnl5Lsof54s8jX5chTM0nG6OSDW9rK0
akdbl5fOviNF6rRj1/OYoLEa+PmHLk+XO+OBN2nuPQ0njDXHvJRQNPa5nS3vfiR6
6EL887NsAyVcv3ZhvmQQHvpZqOWuRTiqdx87Q8gn6C26slQ3OLM47GQ1eMIIi9Dx
q0yNxTdy4dYYXHwdeYbMXE6KDMVcIcUbLW7FZOR3KvWqybZqwaUMS3rAkTG+PF7+
elh6gvE6ns5ZSqGdu96KnTKMfDtHVhobrg3uaOvWcIKk7RySUb/mOl3A9DMlh6U2
tunabfFyOE2zN5fUbPyYYt/F2h6DiF0VSQbj3BaAqfRCO2W3CrsVJ0XGy/M2vpKY
4JA7fELO3yx1m/sTD6ctlYTlu0A+DgtWdduHg8ppNbFWHr7/AN8NtAPemWUCmab0
SnyWeKQWl37ioKu4X8DIj8HTs47P7XZ1r4zsAwGN0C+KJh7FdgrcyLxfHTd2V+h7
51hORT2vDBoqbAtrYxdSs7faOFhlYrOQvhKDatBX8yomZ07E5Furv9YkdAp6l/9c
1CsgG4PXTKGwn+A5v+f1T04S0y4wEhfr6vUifG5iurlGu7jozHGSzK0kIU2CbU/z
Kd15iJBXK/dbiVsZpnl8Bwthyk2Ex9xunFXRh+/JJggKSRXqyC+58DPXJZUjAI5i
JysaQpCm1d6cTYToX5ogNdzwmX+a79uy2HnsR0SmWD+c6PwXZH8wz9AgPNiUcglx
r+XKcbq3WAIUPoKDSxTDP6umdAzndqXecqPx5ICj/EXXQq9XRBkWKSTdeSHuBJ6k
8z0tuPcfnoUJBVWOexbAn36C0A1QEPUldY56UQ+Tn/2tOaQK7MbeECMS1CJVjVmR
//oYo7v9wGRhCkYcU58c/K/OuW72tT1+uUY0GN8VV4C4UxC0Acef1oA8yQwuIiiy
V7J8SXcjH4BU14mtPuyKQDl0+359EWY4I0nRJjAvmJhN/wN8SaL+V9UWYy0aX3h2
W2qhzeTC841rYOn9xIXaN3UXrjmtQ7fNK35erjK2F9ohy4z6hqeMntI7hwFIbLwq
FDsZenSe47Dr5h+FGxp06a+nZ/cRLR0lmoMrLznWS69nf9lX7S+IPYEI7bwN0Uxe
0rqPTokxXDVLSqLqh2JdfZ9mPf1HSJPufz8ImafNPDbvG7BrDOaGYeMf9v3huyiV
sgDK71PRIOaFd2RUpClpPrEs/cZ7XujOjkjvP0Y2vW73p/pGwMS+mhYWrr2XuI04
U+QpFPiXZ4coXtehlZvpMU5tqm8TRTa4NX/26l/bUBCg9tyEZ3xokQOjG//4qt5h
cNxhwSTU9/giidyRxOZHyPv1NoOhV5C8lumvc5qRHNyydVmgrbVTneuXtq32C/Ct
VYqxnDfcw0WSl4kFE0Eii0UxUceYC4N1FwWCF7MiZ456SZmEwLW5QkvhXX8iyCBq
fRQOMPXAeeSBtUZpcDiYVSUeXDccihQDC/miE4RJa1C+s/okRHc2o3tALPVZINEx
xuYiBvWB6WmutqIO0lmzSOwgXsmn5Q/BXbX8FM2/Gn5iobXowvQG6N+z1pikMUsD
iNU9DmM2eeWMxXTjN1a0RPnqhMYy2Xn3XSz/FG0+K7+6nqxGks6OIvYPSSV+Q8ee
5BGP+DevG8D3IDjKgdK5VWcFjL2SBWiOSPRjhf5Awe53JCaJmfLayR5X1dVWYbEx
uQdCHxiJ75quixZu8PJyiQ3kJxxse5gq5uViAVst+qGQtjOD4H8AwUOodmnwopgE
KI89qrDN/hShDsSA9CWHYINS8cWZM7uajxuC4XgydkhSOXUlBG267t/XRk8A3PH7
tNCpj3u4+1H26ak8yteHJ8MGOVSp8fE+nwesD7LkU15vBnvw9cx0k2G5+X5t+419
l1v+Ew1aWzsZRwih2VBlkKoie65VVlxVY9weWZYJXQe8oSGHPDQ+Ep9rNUbEaC5r
XNBFz0jPSHzCuhK1FQBX+k4C9nJCsAShtDg1OE2nJOnY6qrwmzJtY/JmWeoB8vGR
jNMmuBlUIR47AXyGmbAhiBdQiAFQOOQ4CixOyt2l/ZOeuVRPjRqlLYZDGtfYahph
/eks3/QKokDVDrv0hfdwPKv8RKN9lovJpBclhiYB332SSYxEesxedTvLU/XXDSqX
SszlxJuHXlCTIVC9qDdV0Ab12D6CEKsxmfvfn+FLJirrX2LgATXQ40B0myLtX9ZL
ziJCi5cmcO82ZLO8MeKA8N1hpnJ6Y6EE6ogWe1VtoSIvHLhrGVVF3hkq0ek6dH8u
a1/Krccbg0t/9/ImvKIaFOAXw/f5SuAPxTOBQtt9ssLaRPMZyNup6HnH8lKI0juQ
MEQ1AFDD1z4p+U16gAykcVbhy8WwgTfuRSS1UEPgzmlic1lpuDShrFSRC8zKX/Uv
mI5lUwH47ztiMrJ6WV3wgtOgCFsF4i7PpuZ9Htxk5e9m+nlGO57S2GZ69gjFAREH
ig+MnqL6k/g8L7pvXDuoLMJqnE8RK/Xv8165NWuI05YmT3IXacQ2l3oCsxUWY6Xe
eF/mP11RIRi/jPSdZ7v0YhrIXlfNp51vYcRdkiiXXJZJiVqiBAeEZFS6+cxuWXME
4bojLQxlex+xWvSEN9D0MSTB7wEgZyeyB8VyR8ctJ8TgHRtdsGPTrGMsqhgYUGqF
ytx9xHa9Zd32jcR9dp0/5LrOKsLIjyYM2cuvpQ4cQf4OEzOaF/NqmQ0qJKC6ghTp
5qbF+SVtAn14mjUpJ2FrGP6e5d1nXTJDfrixVRCMGF5N5m0ttnEUBdjI+w+ApPVk
ZiPHjwwKS+7xwgiDjoUSVq4zSxrm87bNXMslG+JdcDxslIJIZ6gYykfCwp9r+8fy
xoTyeOYe0HB7f/fYWqd10I1yKMxVJFeWGDtWDp7/9rDdXsed3tBRHH1d5ONdoMV5
KNabZyLygk2qIuvGeNVNvyf+fmmgo6X1LPQM/Xl9i2g455yJXj7uoXugwc2l/SFw
rU3MEmdUXgW9JHCkaOAiBgABSDhjeyhSi7Eqs4xCFZrZuF8YUdhi4wUdpZnDu9v2
pRqeuzByjmqjAuvuDokWFNE8ilQ/irHz9gwFIHp57vej2sQnIW+AFKhIM09F6CKR
adJ73/s7IlRtNgX4Pn3m5vlMbsm98XAW01mJPFudrmX4URoPaiYariW3SYFfiaKT
IAYQ5SdgEStoVSVNMIwsgKcClB/8Fy+7SnhefBRoOL26mUA7FW4aP3nus6+f8sf/
uxOKo3dKbWKxkpEyPL6YFac0iJzlimKwcSFbj0nKDkupM9EpeLL2PsaKCeRHpUQD
ZTe58LvdowIi5yi7J+JzPBdJY0hYxDVjG296UV+bGjXb500w7iIYRP45fJM+0GpX
7reRty0DSoYtJFYTe0x6BRFm3tk4EkoTgntOqdsiBGtzFVS1uUtB8ToBL2jZyxgP
N4DwQGz+vMjvDbJMrCB612O91fvEftSfjMfF43KhCYLfKFy0LzYGG1D2Sczh7HHB
/+tEcFVpyoqtcftzTABA6OPqnoeGMFhlGlrSkr7elqSd6BIk9xDHH8pm7S1XKNZC
0BSzXh3TcrAbA5qKW/pCUgfnJUpL+qM3BD69CVtJJiQ+LzrgOdMn9xyQMO4mw0QM
QgGVqnWGgHWhht/ePe9gm4UkLPrpB1O9MuiaK7KHU3/5Ih9EDKwMhDgsgRrQLWjk
HYLJlH22cz3bJ9A24UxmanfezIjavSy2UgcUGSCClt6UoftcjHPgSZMjxBn/nL2Q
FX5rONm8myUL/KlyYqj1dhd4PJ3ENOM9rEgSTMT+JTptQjlRXiJXowOqIQ1YXAAM
xVcTbwFRNiS65FUaCzz1G6V9+/w/cZ9uSXL6ZoOiK7O5VX9Dz6OoVZ8HIbs0wkL9
YabFc07d4rlzOY4In9C5BEvQL+iCTzO3NaPyXJg7s91dBRvdm60+MFCsfnhsKhgm
gHu4bA405Lgncd7himMDmf7EpmaKmX6o1WzT9td/Uk9XgVkD6yNdnYKw7o0ivQ/4
M1EFgnRkR+s9T6G5UQKp51zPkAxICFwkSpjJkfxJ/6NywYKZJVVOuj81yUHpQQ3b
cDjVJQxeJt8DK+mer3xYzjaoxYRFUCoV3Sd3U6KoCLiBZCQ1WOzmK80q0O8SYaXS
aJa78Gnhh2BpP2x6NPoa9um/dR1X6UsiI3xEUCYWSCMNTXCPm+VOXD+yNUpQH2BU
z1LUf7d1Qs9T6WzoiqC75dmfw9lUFkY9gxnzcmU7rroB/aF26WVAmDwhhE5lpTIR
oOGGT37RHwsopWUXwjCszhWfMDNAz+Ph5xP4HLdze0VsbAU/pnZP/PVVVlb/+Kra
ArwIak9rD2XLGFC3iwhJwDI882yfyTmsUCR6rNln1gA5mICouOnYvreqQOXvqPHQ
PPFE4trhdOoU1gCaf/SdgqkY0HSfj6yDk7Pr2XFx7SSGfHLYS6wd8btseKgwJu60
iRTBU3ergAoiq/ph6tUxUxL7R5Ec/zKPRl1/HpjLraKrJXdTUQCS69R62viIAfGw
hQU1lfYhVm/RSCYIxglkAKakalyAlKvZ/+vDtaw2SAAxGZO1chCGXsxu+F8yZ9sz
bFdUV5V/f8u+80CZDJTFghW3d2E1kko+0Odr/5Pt4tK7CizfpFQ+uveSa4jOJKnp
DylB2vNUxD5mmrlKxfRaddPrcTuRMItPE04rf4xnw+IZQSihc3A7ntCeZ/Rlnxm4
+t5lASjHFPVvlgvBSyNBsZefdi5zLjfR4apQjJ60b/MEcLiGUihEh3BncNn6SabJ
dNWkcS0jWyHdWOXqS4KIrdVrBTat/8mnK2xtZkoilxe7mS/HC6bULELzF+QuM4fJ
A63IvdFeNCAjqj1kHtuKAsB7iqNx/bAkaqXMqnSAOrKl1td69hlytCftvDmclxuS
GhXit7dmNPu1E/AtPzpa5rT1Z8cf8X5/GNAvJO9JXQ3GKI957ZdG2HR1KthuA3y6
11u88z4Z53fyf+my4rMJvKQntDBqgxYieHo0QXHrD8h3Bg0ytAOOa1LkQqyT2xjX
AJ/9VImTWruFggh1sge58N8ig2E9eLa6Evjdm6b0uln15EkSfZ315EwnB3aNHjqO
8teBn2FI5eNRcx0LH/KLPvHLa2CfpqodN6jFGfhijTh6zylgJtkyMzyJcO/fqeew
Wc0nOrbFDNlBn3d4BPyh6K39cVloOjMbHx4PKLOJu4EMQKoeWHbQjqX3pSV0Ayfw
7pxEtVqh01Yevo0IHwvv3Fn0uBW/8jumloNOClSxtGVzfGn6xHA2tfDUM+yvTQev
EiibKuvuHz9/B3sfIFxyLj2cG/Dwh5X/GcK3nLbjQCuIacheURpHOylB+Yo4I6YP
+8YsGtw1xQ2IKI4fFTGWVCx6yEmtWhKNsb0wsG1kBH51MCgJg/Fj2pxckGOzLdVe
UQzP5rFj3yQ2NLvpOQNBB4CZIZpWB5JtZf2wwUCskQhWglR9drbRcTR/EcmYxgoD
g3Umw6SExUwc2kdLb8EijwVKv4yfRLzCjDCeWGT2G4bE+mrI3v+4/wwefjL0elSx
xiS9ZOhixz6SLeo0gaqeknc+QdTq1zsqNBcSJD1jxfcNOWeEgab1IYVBmozbxVfW
E+5xcBGiIWS/4bC/Zln/FbNxim+hFegiZqGKgrTL3IMjy9iZ0PTAzb/ArIaJb+gQ
OsEU0P+gFtfroY4MuR45+7WUHsWXMlTgvItz1DtTdankQdcuKU3U/izbsPVHlaKg
Zq3vepvEJMDCarmLaThlhcr9F/wxFWI7KjK256CLBZZvg7QUrGzp6JcEf/VAY/HC
wi3NZjVJ2LyqK9itOaFNl8U7z8UkLRuqqisOAk699tXCdt/fr79NDbA4a9IwIY2j
DYt1v6mj8iyaZ3x3/7HCGh0pn+jmSKcfacvBYZH6t11v/FFkIqlKO4LnIAY2kKvB
AsCGfbmgUnpGFfBURA6Y4KQBe4k4KG6JfVIlDWekvHhw9xq5Xlkz5lu7b/OQkzj2
N0Ov5CjvBfM9ASioNrdkrgfmG5xXHAQ/0ToF/BnerpD8B+72q/iBqTm/lEDjSBXr
ZI7inzITNXRFbFMdxZ/tuQhNxKzMntCSwdBkTJYbDb+QeExuUPKdKyQLBLvxuG99
yitx4TOSupHQbFzGODWttuLZCuyX6BsfZdbqehxf5kUNrLU1OCy59xEQToSHu9TB
1OH4tNLxz64v+PcEjtESI/bKchLawhDoDx05JCaedjMHmojad1yD2QgbP9j3r2hk
vRGa9uP9jxpzSWN6FAjZfj+i55OWRKGeS5HGCye61dy/uaA79j/RUDKvdhEV4nNt
CeBWYlTPa3Kzw/G05I3rvMKFowNaEMhIoNVeDmAHpNGTFDxww9OGo7RPxScd8Ljo
r+A7OfOY1xYGAWoW5FqGv/lsHbs6X7t2jjS5ZhS1K2z91K91CF4fRy75YlXhGAFl
6EBXpoKNsDFjI2KWXIkxpE8YaVlDF1LXmv37gqFBrdKTvgkJca9BmliJMqnvu0ib
ygbabZa7EUPGNpPfNDwpJE2edMbXgN0EiTJf42clc+7lGXVubGxzxfSszAPRqnBs
T7rIxWJ/f/281OpGB4oDHDd14XzQX82dVhx2DoAmY234c18pHHuhAyaNCMlwZDkm
fpIph9Ee9R8p0Q8N+3mOmT6tragY169SvHNMauk7/ZXznOtugRHiik/XXzU79k3D
tN3BS+3QkVjmQHcI2sVjCjaX+jeTBAJmhNsidexHYAQIXavbJqIDI5aYfLC2p+Ao
TqCwatFTuIs5DL8/1Eiop+N423W9l+Maj0upWzLwDKc4moJaP2pazgFj5o/fDmsb
V1zvG8C+E+8DnCL5gqA2epODUyN+A+yl4iZ4FuOF1UJfbesE5wTfAInAYT+karmo
tyu92JPy47dG81ybgwDoagKQ+h0Y16s65VVVw6EhATKF9o4UhB/Zr2bv+qvGLgS+
Y88zsWAgIXFZmNZxOEbMDFVFqt2Ejxx2r9bfI+WFZ9xxoAcuo5HHjuMYzDdBP6TL
FOMsWdyRHj61Xqtf/ZWyyl96V4N8ucZVvBwW7UC5lKtVKS7zTEps9zrYygoX/CgF
Vd706FnaY5+IZp50nuk8nVxvMmUr4f4WVeCJnF5k9yyu1j2xsFsTyQGvbJs4H1Rn
ktdS4KVhAuqWyVfbEtxoXxsnnQFVjlM0ISy82exuCAzwgCTw7Cer9te1AH0lmsu2
dTWjCbiFFai5wDcObcZHC1hIAUST1sraEMZ6ry9OtHHMV+Fm/5AQUITWP1jy3FIe
no+ONoIEArovtOFK6uSB//zBj89lKYQElJ3yIv18A+S0hP8T5r28CGLwZoeJj4TR
azGhbSdTazc4Hj6nlfH8BFzGk+OdhxUuCC93Jn2/Ka/Jz+zJlZ2G64kTCZG8fuwr
1CIUBe3fePTHnRH4b5FdPQSYG6X0MwDhrb/iDKU4bwPgYPNRIS66b7cV/cMB9eDa
twIC5Gvhh0Qyb/o/mvaIKhsLtnhI+DHpcx+o4OcUzupRQou+Jz+7f5ogYhJeWgXz
dlXLN901ODULcXIj6lI8pyPxvfwc1HokrIBgDjz0A606hfLeOm+QB+HdcR7TcAyE
d37VNDNxiSRj4rtfIi4tH+laBa5Z/VfLg46u2u5hwdWuQh5uoEqR1Y44s1l1cfi0
wHoNEkJDOOtX7vnOfgDwIrXu5jYRrx1kbFsSCFpMhIpK0y5yQ8FCEToamEVIqbJU
FPWW5dzH8sRn6eFGZ3wJXkTRFOpv2vr2+FbsN+x6Y4gV0cqQ4zXzVBvppfAmb4fi
iqSJlshDEa2ZA09wFndHe8h14zzFMBnJ0YbFyYMar9zZsnw79F6BruxFA4XDf+/3
GGxxEu5kj1UXa+NttJzJmNEtYmrXPEARY/tOS+OW5hMYJEXQ1D4hPVKuukQWt5Sv
trOajRNup9TgjGnBgKuebmsQFF9+iGB/56dAAJ261dTXg27YOba3VRkJJwDp7N8D
ZWKgLGwFsRBO0Pfm71glYeqW29u80jB1mwH+4m4bfSb2soW+KpoS2Kp8ZdUKUq9S
8akfHzRgDj9jm+lQuAXOY6WuJwwFXWjXTbV3bNntewq+j2T7cTgtHVzFT5xKJgZE
7URZboGgsfowCweUJC8VcO/LoMwDhOHHOebH5YKez+jyQ0dbGETL4kW0U7b0aj0+
NCG5EGah9g6RAo2nVifLc7JHJxJj+YE/ltSK62gSddFO8zi00QVKZhO802jNZkoP
Kbui/TvzriUywtwpC2rOaCgJrgf4r7RTCHoIzDlVd2NBRQdG27ALrGG6PZBZ3EmS
XchKAwwxPw3F2VqKKyluuuOXM2VPlMdwws5LGZi9AG+BCyig6jKNeqYBYV3AE7k+
ILxqJfbA2gy8gwx4r43BRQ3n3sCtJvItE3hYoXLYuVUTW2FBwcBrzx9hlU7YyK+n
IJAd3IgxLdsWRY50ME7aQkqGA4fpMaIfcUEXdvD9JfO3bn0++gMfj4MWGQavYrqA
4KkCjzbVCCQZGnvdb2cmovqwA+rF9f3GefcBsMcRCoX6gmjyrUYPxSNIfhT04JT3
erL9NZCKHNvFOb22PpmUugIzhSTcSFMowDdUR4thfwW3XVjMzd9Bdsvpk8YQ+R+1
D6KeD4s3CuKIUoO4PaoSblFJvWJCEQl976h60l1+mdLMV5UnHZouxQht+VgNh9LT
hSiCDSSURRfiXQPKtGN4C8fPzLsWwlr3RA4F7yacBrPQcIPIu+dd9Y+pIJkG6Dev
QTdGCKiAzKL0Hsuivs9WJEY97mmkCJ5f/r01lFvh1o9qyJnRP1ylZ8y7dG5TrBT0
NH2FFgUiAasWesEB0f+suM2n8SwRnKZ+VRBFKyxCT/Wp0u/Ucl9OyFmeNUdGxOWx
9OJTYnHUQGu+fVOkvjsvSKZMSskLchKEp0YdgXJSCN5DmmngcZiYVKHhqrEU0VWW
9ijRTPgyXarFxQ1y7f+iZPK78rlckh7vlKCSfEzYbkmwMUVEHo06+3rnQv5xfH/3
DSqAOLBukpG7lfsr7iqhcYh1gmLW2pfhUQy/3YL1FTkHxwDCEwcixBVK+wFt5oQz
1qJrJYuQlY/FlkliuPeNJCCXhQ8T0UPX5g7vtsHiiBlKQC5abF0/Lv+EWdo4jN5V
32bRRNqsqOjLTYoxUIcU585TMwxnFv7N7TAcgvTtztjcW5ydDUS9XN+VsOXZ9rn4
bdbUviOg5facNE8opLebDBZeUJCsB7cHxd5Z0Xe50ViQNuPyH/w2NVVeD0wi0JW/
GzS2dFaCln3/qkkRFEsvn7bIBl5+GeoGmLDclepPg3x6ysWsiNdJpX0k2mjazsL2
eRIp6nuveRxUmn9H/Z4Ttmx9HHa4mxGd0EUVR1OIdhI1q58QSRuTcu8GHtZUghAu
thUBEjcxjc5/SAlgtPnwdhLArIwJtLdgPI4saUlPe0HK6XMEo8kUUW7l+nvATjuU
2kCcwcmD7UT8y/RTceqC0dSl+plSvqHRxeT5bYzzUY4j0ksOx9qrGk2gvT90vr0o
etvdW4sqQR4zw6SqUSold+FLMNsn8jZ3nFHcnAwSJBblUfqXivTe0c3LpAjMDZJM
+hiMKNRfg3E7IgFdWPdnKw5bujWxeI3iNNCwitABlmEkxr8aBviNuyOWSx40K6wJ
M+o76o8ysZN5qmcsgJmRyItvYKFJZBdqZyAWP8xk2axsJm9FKKnIy+z6t3itnHBS
EJXpQ9/eymCPkNiNYcZiFHzK7JBAGTR6htx6OChepqoywRKMBSCXgcsgT56T4aRm
NZiKtQ3N7q9GjU7dGYH6AhOjghM6wtvTbPgH/Xjc0OWYgQ0EdiORRkRFdoaSgBBr
bCiQxP0x/7mBQgg8J7mM32ZiDVBDFa/LBkcSIHPTxPNXjRTM+kkjC+uoLYIt2vMA
H6TKVRbd+Inkv1xbxg8Uhu2f0Ow6jS+ywan75JnSUSmCx2XoZYQjhZ5jx2CqQ7zF
yq/2gp5r4vTt6j65uYn29PEI6vRTovU3i8HyfwBrZkV2s4uRE7gZhCj5io7QO7j/
pa0swcnFyF0pRRcydFpnZEMLbHU+NyXxP2MO/rYs1Rvy4cDukveaILgge+I0jX0Y
tec4E+8gAg8rJ9XHSvQVJd3NInJUVx+H/1O4q6v3usw8ZoM8HABygQtXWWl/6+NX
GQUhkXpLyXaosii4oyxgmNiGT7Pve3kXXzV74nu438QZeHYVVAoqI6b6wjZcdHRg
x8Q0RfmyvA950q8/JoRAtmj0mQKdBO0ku1glKJr3GUAFp6lEBN8NCdajnS4sV+QG
QM8jelFSWB1Y/XnlkoBL7/oqAJiKl99BKL7DO1KpwpvkZwkI9EH0IQGuk+/MZBJu
ykIWX7lFTezdMndyfEXN8WF6aG5hTEX4evRRV04b9SUARco+mGnxCHTTy03+cMpT
tuiebYji4IdI85c2JuOsAnqf9Su8B3F1qz1L4hj9VPvCgy75WtQfQAD4XcmFjpjf
vwLnV54Kh+hClaG5XWmbVnxatQcbQDTTC/XSckrTZh7VcVpBwFwOZPHi839zsssC
q5Y+8u19frqt9ZKUuW5ShlsVigw2x35tjyieE4hKZqJN/xQJvw/MuI5tXo6YRin1
183oSWSVO1mCOm17pFZO1OV9CjgtdzWObPkobdhYldeMz1rswBHl6d8g/WDzoXLs
/DlLIr7ALbyefHbDUKa3eeTS4r5HYQwZUm4j9Eeb9FHIWAyOMMTZPkhPlQk014DL
mwU3qGNYepezLEo6QiPuwPdbDY/v0ODhx0HmaoEnO8qSfqQZ9Bw+kZByaExfkQRP
HZ2ws4K/jgjFhIoiPdMpmcevYFWETLMpHpMDBeWAa5Jg1VgXlTBlA+4kVgm0JvOq
ZFqI6XAyPlQhGUZ0Ztv3rmikweTET/qzf/V891sGXj+a1/hWwpfnjkisZXVs/qjF
s45ApUzLcle9RhP46iofmH17toY5ZA+J2fx1sPUcqsnNpZTshj5bmWgTCGIRdZEF
UkoYryZbZICaxV08Qv6hNPrncu799aPOvMlS93o04jbVhju5jeggyu7mBOXlUXhS
ytwD8fiAOUEXzShmru+Cw/npn5Vta56cEwXC17myEgsInW2Leo9E3Mlaqmz9ziXd
P6cw5ED8SR2Ys8v28WJdGfAeb1gdi9N3K9xEGlwpAO5fzwtogQY8zfGf81WFofrH
r6XRHd4Se372j5HvDel6NEPi5RnPFX9HA7C7XHq+0c4Lv2pcnGbs/s3cG/HeC8K4
kaKKK7uNpdTc1jkYJGdZStfadtzl6yGIjfseeDSps6gI2ygJsgro6VL7/Hf4bfJe
q3KSWJHvUZfOqTYt/KNX0mACSdcBkHRqPBl5sSP3efleIstia4/rerkJMiVbWhIN
47aoyhZr3tcIVCtVxL50eqE1e1Ll1M5ufxkUgo8JaT/IiYnk+UZtEggWPxw/Heyw
k4h3XfTdHI27tEuQkOt92c8NnxV1BQU6M0jPcg7bfDfywTBGptUxdVU4VLugDRO0
l4qpgi9mTeqrj3wBBKKBbPH4myU8Z6uVVF6sfUEkp9PqxKhJnvv2LqXyw+KIePnI
hofMfFD50d4eo0yc1mzveFZztQuIeUpAY/rN+0222XJO1IYXtF/S4GEDfnmVnxnC
NwVNnc9/GZdDGe89C7MRpBp+o0BZ7A78HraAbNzszGdrcQVDrDfgqv8zxz8sVuYI
7CURwrx6qFCSzlIsVgy58pcQED2cs43Fw2MHlFOQ3O/13JMBSGSpUcXAGTU/yivj
7a2Iy5+fbhPjX7FUUxg9a4Jla4deTErLw749y1dKYwHfdFA+mVZubrIxSFJMY+QQ
JCBzmPTpyWpE3M954YHHeNhYPBREsOmKZSHkrR4g7P6DPz5RPyMrn4MDCIVL/DSZ
Bhija8iDdYWDYuQyilyJVJIiNeTj0qrODqO+ZJSOUzUDyfC8sQGgVlaMMGh2BR0Y
S3zOKTVEEP53Rwpzp9CDIF+2NBC/6sLfakHmlBTnEzcNpnjEGo8HO718pZl6Efxo
K+DmMcmB0y2gHpFxzN5wsbtdGmctqogsXzOZNhZpNLhdcBF62msVQIYM52y4un0s
UDF8oTvlTddNhHBRmVncDYHTuc+DbJLuW/RH2h+A10bQY6iKfpPxh0Lvld8n3kPZ
dNWAWooWvCkQ0EsvH5WnnO0O5akOdB4g/MTW1BwXlvUXsdNSnxV8E8kYjAGhw12+
oy9CupHaeUu9TdZOo5/dGyI3J0DpUumVyAzccCqHm6t6hU+mCyRHzzLRi8PD++Pj
Oa07RBfpv7u5Y7QJQssJQJIRbG5sl/M/jXQz5Ok7LdHyICapmOQ0VG6Qs3qPFlOV
8AtJKff27fd+iB704dxgmMPPXa499o36XvpYGSC3vXclwZyPQXfMj4DPNVHi7Kqs
hNXd03t13M/oVKG3AdoN5PXwH/nNHlVpKnhM/uaw0XfrBdwkoLYCf5mWavGWG7qg
ok7s318uOhpHSQxyprdHAf0vqaC1lCVL4VWW8v2uUABPR8XzmNqIsotHo60N+E1L
WC29LphAikPgq6u36AxTA2b8TNnQF21iz01wNrsa9NcG5G1qt3IH3MLzfFejfclt
DmFUwGayMWdBGS7gzFmkDJRRtq84gBVQXVsN3kdoTmuC345zs/wAR1i4bfVVhUNr
3pun89SCgzZdEeGoV/TYNf4mJ1zWtX8uzmO/OwANMKKsjckMsAiBoo80D97I8QQW
SarMK6Z5MVl93jUAcQ9d0ChuE3S4z1Dy/L/Q+MvRQ9htA+NYdyj0aXvQ43azutzx
PjFTLGTUaqclmmSdt+VbselOICb3K+eAgQsww5FASZUwM6qEPW9c+gq9wzA5H299
GpjCaNPXEx6vw85egp4FyRQVTnbcPMJ+7TCZAongSMMetNHtuQRqXqeE8dUKiWHA
/v+LGg9HGdnP/Jw7Gc44I41pvCe8tiqWFK796wWR4SaUUVqmAbJ7yxumUNQu1Ysf
G0BWqNMhhLnW2HoudKBFFMKzzpMQwgBAZ14ACd6wbxfm/4D98blZh6gyU41/vMxC
m10xPx4JfOc+1v9H26MJ0Am/hV7iFZUOZGodpqafs/u6emFwr3p1gViKue6ScqbD
8UrhpUSrgzMgI9oSqEhJ0UWjqe1tshP8fofH0j3rqwLefbM6ckHNj5pH1ORWQwpy
LM5Lvlb14P3/H8hDz3vDseENVur+kURFd1FNu0K7798GeO3Xw3R9NsdTN9NKE5IQ
ABEmbufDzPcUtm2XuDXu1wSRXi4JTy3YzwyvHLgxNVSI4waRczzhBeQjxCmn4Aek
DFKnEEaDjEN5T2fHT5ML7YS96khAUIEtgq/kBDp6wMkk97mpXfEtOIFozKDYQkBc
Bdmv5zS/oLsggtU9qHU9mTS9HvdzJHhbkTtkvjsnBUMGqNVXDvbyMIlXDh3E0VC0
HERr26qHCvSdR62g4wVaGvAE91JWkLZNrUfQ2B9IIYxKfJdDRaJdh/RQuzrW1QAo
I28TQwT6j7fo/AzLzfAfgcuBtCkLxY4IubHcp+uEMrlAbY4a9fy6hcnLnxbQjGYN
l/AkpUtTGWfq4M1XUquWaY+o/JK9JJ2TMZyOsJJauD+eHTNQKN1/YrHXdkfrymr1
zUpY0W9tTEkr2K0ILDSOYgYAw1akRobVv7sxan/Da1WtZQHNyIKOOJ1L+CINMHvg
9unWZXHgiRucVr0khYNemkNxE79UQQry26tRlqNO6K6PlCltUgaLr0AIR8PVhmWN
u2NhR9CKleYhZksqSTuUXqdgoGqda/D/9GbBByEYVPX1nphKiodLkv76PWEHI0qH
7JXuGficbxerSxO4NzqLBlVOXgZK8zz0LOHTUE8Vu0tsPq+AbJbhTMc2I0efhW0w
jt4z0sVD5WaYXInWuENAyhGYXfUP/M8sXC5WVH9fikyUvjgPdHDPuRHE9sN4E7AM
6tmMSSatJMTnO2feFTpkoaHytOvK041bhQ5EEd+EKbj7wctR+X5H+mapFLkCsO+u
0a8pwJ9apCPOakDswCFgEy0bedQ/yysB8QwtAIt7I4lkwUsZ9Ooo6nEDll+Pdk4P
9OR7UvzVEpzT6o5Ro7pCuJk2DbT0XTDaIT4wIfHRX0l8+jsnmrAtfHGxApKPuug/
sxqZVZcZmVcRsLg+xiOlvlWXhYsO8AtH0iqbBs/ploWBnLar0sVPqSG4M3+sihHx
5QYESdA+BKEbbif3j9m+U8Cum3arH2kLGz6FJO3VcbwOQwxpJegyGRTSadULD6Jg
P1Wtb3UoBHj2OWDlAH3OIdX0xhH13WnRF1jHboYgoN/32j0T1vyxdw+6a7jd8kXf
+DQTIIpKL6NYUCwolXyVs5+hXVstbrls8BxA90IReG5XFU92/m6pW4LZsiwxDDzj
xCXugkNEHPgteCGLStq0DcujxqfUwl26DZ8YSSVlJTH+Su0xa5gYmvkUGg0yDe4l
ab6LAAC5E5h4nUY0Jisn5kZdcrK3Ow9/d5iXFkCwjyYH7xV3BFhnjYZgxV7bEqFa
lMnJzzUWd3Mmr2aiE++z1IWYSpQ2MTIPb+ebKeTEaLGRQJwayl7Y3qyuG1hXFa1Y
f+GCEg7IAdt4EC5yQu5SVwtJ6qXCk895PnFb43VByaWEHaCWx/qh4Cl9QXxGjG1i
yFOuxXP477HEXa1jL3cnIHfsK9jn6VDScpLDNYFk0wl4C5m8LiYuPWf2Qq4x6v46
0kjmBYJkXHsCV5pTHTHKURbn60N4JdkWjkdeQtss86ciiro4aXkp6OdvPE0Ptmrb
nb7gU2S8C3vkVqAbGSgsZOzmB5xzg4awm3xj1tt5AtP01N6xgUSrnEZfCtVUw9qr
BvkKhXdMhokeSiGMM1pskJ9MT9lzhJuP0YqleEqVaWLsAbdEZNnwPYa37ATXmJBH
P3PGNwzOvs+3zpIz5kzAfjSE7k44/pwE6icTpF85PiElyfseca0CUKPo8L3hy+Ua
MlfnkWMfjeVGANA+8QHcyXbf3aqfZCmn/e+a12iwmiuCJC45s0PCw5PN0nz1QZFQ
Tn+3XbsGu5Z52BCaulnKPzbyrbKDlBdTUyL6pciVydbn9jnqe9/2SuvqOJaey5fk
/WHjCN0SZBf4qeRre7w4cTlZHxJqA8+FFMYnvUbB3bHZheXi9gz0s+9GUmi/2+9j
bPgl8i4wMfX1iXULcWkDjVKpgD0WNIhXM9m4KNpAp+pMTgKZJkn6vBB5M0FfuHt/
go9VKJ+Pza8Xm5p+27/uqPvEKCNxW2AWW4M1ZblTtbmWhVO/Q9V9Tk9RZJMn1SX7
ewnMsr6g3wKTNia+l0JPl3xpGrSbffF/7us7Sh2MutT36Buw5o3PXyZ/QYnLSzuA
bwVI/4dNk86+GsKPbBYRmVrkbbGWPo6BiEEASygq31ju9/6EqLv/6Q5LmrmSYBxG
4Y5JcrR8dW8T7k/FbLZnPD4clxU7PlBuwZRDKDFNaKpD9oAzKvmP14LsI3iQ4WBr
xqOoHNuIItyWrYRs9fs3g88EkLvVxEMBfFhQaGuocqBeiNjNRiOZNWAAfrGh7Bd1
Qj6qyHLdI1L3gF2PKCtcLywyXtilovhucEp0x8hW6x05X1HbFEqif2Ug8I6NqP5F
FuIwabofg6hGOq3af7pab2knb5D2e5QuvWdMeHLuSE9EEk23psg/F/u/FGwrfBQS
ESdmusejCQio2wC6IzkOxn8qFePyCE92a6v/dv7gSZ4H688ZLJhdYpDCcQ1YBxlr
tjtjp6UZtz+N0Ad7rbYiHAV+j7afQ88ykmk8AakS4JJ8DKdaE6clnVlUbadfXA0g
PgKQoxqL4dF0wlxUVc4W5+eWGJJnYFtLQ7xUy8XSYdZNPmx6OQUWDoZ73CVEBC5Y
hH1g/RruF+eK3hebHF94beD0S7q981tO2i4kQms4GRmQI39nsKZZ5SVu1zbjImiE
rnlPn84so4NT63i/Vq5AzY3CULdqe8dm4bYSp+XljXR1dVHCKX1mqIOTKRyYFNTC
Kv81NToMGVF4/ntnxBO/IjAs1lYnNTYtttM2+uNynx4+wdhM/YsEEvYKF2xmGcxN
Of7GLb2DPugr3/hb5n5DN4tPEy7ai/URg6XA+Oig5v5BJiBaxbnVqonE8IuCbJid
eNHwNoeylOgGJTWhNxDhT016CLtpM+OO8c268os4Mz/oAvbGWOJh10drm2X72Eax
y8h8UFA3KY1s0MU/rL1RGvLFITp3T8radnE9BBri2FIFaY1ANpgZCA7eA/2jztpq
Oma/na0bsveghOCTwpIrbB+pOw9XtHyRhTOnVIkkmSXSUizd/MQ2O7+AJ85FVP1c
hhqf3qwrrBjWkXJchE7KPet4D3nk5agPSWKWtM3Y2lUHJA7dYc+Xw9dHWnF4/P1v
rCsbnxz2f0Lr8C2iOzvsEHPXqAzA+9QymzuhCZPgZOz/3LWoe6POsdLPgbHAAwJ+
l2TjBjn38dg9M9wb8luAbocesLZwPtfupMD04LwoUH/cTuIWkzRcmv9lhwQIMUC2
vBUST+AaTbQ60z7rQn4xEFmK7LgLIhWrhVYgb6wr7a6s8/a9NyewaZjFtlaiPV2U
Ep8C5u+wBMw+3Cq/lYPEZXHXRWcOrR6/jEZqnUTuSysXNMMyofjM4aH0zUkw911O
spcDXu6zfjCRH8Nw2H5seZmoaYlU7WSeJmCzODRYM7p7WWt3LrSRDznjNeVYAnjO
/+qPzWe1FEsDvKSZDomw7Um3n3cHOFfc1Fzz4zLJqfmW2zPOfgNglIq6BCkX2KT6
kMLh71AgHTD2/O8uEIktuNjXM84WGE0g6UCdMhb9Gz7Wi//TgeJCoEcrhS5sEY7z
F2DPIWkvCgxJAiigfcq61GkHEf+DzMWLXPRCgzLGQqDK1krYtLVFhk4H/tE0XICL
gFI1e7TEdhAMVMBe4IQBu1QcX3bZD0He3NQNiw8CKnd++B0UGBGKCQ6+iiCS75Mz
f7HLlnZqpz08DqqrmKYfzUTwuP79IgC33sUR79jIv0TllZdbfxCOZpOUY+cNIqBA
3SDTPWGEib+LBURz9FUU/j6Z9RMECc5regebkpJCOtassiJFKBTcg0EcPjaQMDDY
ePBwaedjyBHdfrtuVNghkkgzZcZp0GoxPFvn6tm+iv/fO38uIOzYG4xGY+3fYFzh
MVMiooYLhkzAcvEAtHNZg5K0BR97oKgtg2LgGuonG7bHrkO0UvfLwGKYFiHXMzde
2afadF88a416NRzEkLWSNviwxSphgXCOvQnHWgTMYss+e5InT0BrgFsY1R1AkZ4i
IzGMdFyUCR+cpKk+pV/1GBFiGlbaTcKbbi+8nUrw9ARl0/xtC4PA7sfGtxhnfdWY
hUIGOfwvcu5P21dDuCh3w3e2wKkFYJPKdgTitISrP7ZTPaA8n97HVtJd3DGVY+CZ
BudLjiLhqRqfwtmyjNz8b4baUU0MlCOlvT0Y+78Q0vaAW+p7v1ygYC1ffviUHon/
a3FhNpe7K/3fuuKpY9gM433htYKQa4VC46yjEKHc7bdu0EZ9cwzD681vjlNPHlZA
Fz1z9dRpG9ZbNnssAXlexZbqQ6iSMDwR1Qez1QdHDczxTO6/aU3ktstKsWgi7gSn
5QuT6mcazb7eCGJb5fscN/ab2wBbT7noF8zArvY7VbZuDvJUmtUyYwV7Pk7ovN+5
6GbBtqg3VgWkqEIuBIqb7HRPiayx5Bim/HneF95LLf483FEVBqOwDUVgB7I8/yBs
7zc7aWhlIjvuEAAFZjjgGbl6a5bZMxQzrWT2ghpnhrFbfSsYQcTXOT0n9O691f0d
/sOYotQai+pWeFpNR5tMCgsf3474d6obJ+VPY598o5kRAEjcmAZalMwuYoPd58j/
5dPxdgkIBcewlXkIzHWRrz6fQxP64gfl2OAAzHHmFnSLaMbxcCOfxXS+Mmnuddlh
cGgnkx9m9JX5lEOeCv1IccTl4LsIzTfVg0D3nUWx9S4eHkO8kSSjkFhziHVcJpOA
peyj3+M77hG2nJaw1SJuHEKo2NIJrH9xE5tK2DJCNTDnFhuy1gikcnLHoYk9D3rR
p2oYqzuKYg6fiZrgNWIxk44SKArT+ItLv9IkTBcFJbrajojmlfA5eEYW+WPwqxTi
fT0yBW5d7eEymPpp88ENAoNOSdKMkc8DYp4FlqVI8XL6nIbJf4Axs7Ib8rSfwaUu
d4X84VSeZEQOoTGqlXSgkCA3C8hF3gZtobCzZLD0ETfr1R+gMMJAuT9XkIEQb6bZ
5Qe0E96kTpowSICYONcLiU10lw3JGe0kuEXmD0vv/fftkgqhu/cvXMNbJWd7YoJo
ouZFA6WneQiFyprKf4pijZeSNC3cH79uaPSWOSW0H9xykd7OMf8aCIpuWWP+JMBU
cCtwNYT8sZZ4qX26z/SO/IanqaSJVPKt6ilBaQrKjWxiuHTzcoldXQP3VP5Fye5X
hZDKqtts3WTL3Ls9xC/Nj87wJ/Wkv18gLyueY7VpV7JxESflA03wnz4sXCxwu+Z4
iMyS4h0RtrstpXKEWBGyOGm5GJIeXfPNQmltuNaIaw+Sq2sX2lDMbTlhBAhmt1it
axOIRgmLwvGFxDhJpppJvCk5Dpa6Wm5Y1CoBwP3tOwCLGfd0+Klm4Y2iC+RZUl4D
1x8hKZRINJuLCdAVqfCcgDZ2T3aEIvRdpFcJAN8ahSk354Gico6TBacS/D/b2856
gly62X2Ty2TlrlPYG4Yai1urPzzK1kQpajGkK33Br+VFXoLZmpcJZnJpZtYBvsV0
O3h1i4dIjGGhqiGhj8NSaBL8nQvx+yT2Eu9DBtXN6PnI3MLKit1qiIiTKlqDVRYr
P1gMlkBaceu0cKM3bz+k/JwuJA/88sudKttvt7EQFBroboS29CAeDuCPkTwXOoNZ
9ankRAxwQFIruGpyBb2w2+lXH1CgNSVBRmXswUxnN6byBpaMza8QYn20xqbQHOW/
gk1WZt8bfjikZVvfo9jnREd2epTtbCe1ZBxrWA6Ulf88km11dGEbeVKqyn3NAFlL
dwsPbyOvYz32IMiZJpy2owSZwlYTo1c+dLQX/HA6U0Fp80fszFfb0rPR7DJ0ogxT
cXNLNDEPF0dm6+cEc2ITSiuAFJO9Oqr47isQ/sYRdFbGTjqEmaQXoBw9vVsHFKAJ
/cVF+aJ6ciIMyL3WntI+3gBdeLyWTqW74JZWfDL/6YgtF5f2Hz9oX0rr4/KNAe9h
HFe3nLTTS2qTtZIbyQHeppYEaR/lZwWn4sKSzuiv/Ot/BHHQWN3CE1hYbsjbAirJ
NwzG5wIgNlRUT/jP/jheqYBKSFaiLSoAuo5/R2hqY6dVHAJIaXk6yolA+DorkZJN
BydIFGsF2/AVaJtEjk2ZAcH/i8oLXy4nwWcV6MMpEbCr4sygb6uESHWo6zN639pS
ljjpM1k2n1Knkb2skmjKVSIkfvh6I3OsnDikln5JFbR/UNndxavCTS2SJWs+1NF3
ldYPneRrGK4iwrTbnaZVyLg+l95FTVFfrGltoLL5EZSwdBObuDc+cnC/SnsY+JVy
dt8v0QvD1vfeOidBizg54TzQN3AEeYyn6Ggq3x3iJ67y1HueeH5tOtWcFdHqwOvB
q3kWsacqY9dDv1siQLD9tAUcRKA4JtlAzEXQ0aKrkyNebE5hO1HcHTRCrHV7PQ+t
JS3Fb5/iXzqlYaUV4mBIBqxiaAtFDej1lf+BU5/3cs+8w0xSisLgVMnDsMoLmAST
dLsMYnSt5rJ7chzv/2eaL2VlYZc92azscieTqm1jCKvzv3IwOaMIDu2h4bGB/V3Y
hPpJEtLoCOPpHqSPN1F24P2nOy0HGU0GNKeF4GVvpngPOnxxc5yKDHddIJJ4X9ls
nohSV3tKGLJVwCfegftg0G5ccqz0yteBvxMWk0xOeIJE/45bpKuAgCQh/ex4aPe6
ust9z+wkvlIf40o1djwm9aVoohkYvB6AXAbKwWA6RdpoZnLq1Z9h7HD1KSxUMoOb
7iAuK9/hADbH3pyJLrfgWtjEv3P4SuiR1Ii1rE+hdcggJ18R+9YvD7BIAuUo7eh9
1FW+vT9vX6gutYSG2BUbNJTNK7LZPbT4Evp7fLfwawnHgi1dxfuAWXYdD0I2J2hk
JNkpeTez0+f6vpn+ZdjA4qpkoKXBc4ky29pw9y5G6vj0BHFJNX7HPwB0UFVQl7mt
xORv3V+ge0I0wWTKwQX1r/IO4fWgR8vcvVGe//Xf1hpXRa+WsgCyklOTDpWDh0pb
VkuoIqHGtRla8JvI4SWIycaDfIVvubB67Vx/GpVM7Uz1oZa/X7iX+uQuYVY1a4YF
BznSSVH2Yg4auEyKJqCtHUKdMK0ykdpL376ZWmHwIjHjJYCAv7ErjlYQew1WAgi9
IreHmhm7axI6b7LNOqMezw0GqvD+O0BEKB/uB+X4qIHJE5C05Lv/jduN1TqFzQ+a
ne8jmKO39GUg817Y7GAklW0Z8AbCjIjv+dtVzNSTsveTzITPLsqMkED/7kt7kM3A
wtASAWyJtjmQReZUZzfR88M4ALKoo8W7e2WNp8IZNGNLB8WGgTcFK1j1U/oCTU0w
lrv1Dp1xKgll4R7gj/sqGBOe8czQZIsQT/yitEhPiT2YJw/tt8mfwPumN08LCwM3
/861e9k5bCVFA6XMOZaI8MscA+Cp5tqmhIiAC+JF6zWAs7IhFGdeIIXw9ApzMnyW
6OLnBEWtd+2EbhdWhy/WTS7M8gnt43YrW86VISa4Hr9ifOZEWYdXFbD2G3F+XfMD
rCVKOyrSqnOuA55x9RE1NCmlTHlLckwLmkRYdp3u7DQa9Hg9+vddr1GaO0MfeL+7
x2o2pifM3xRD4Aq6tk6mOhI3SSL9eWPFPCpAEEfXhbYroATyUD/YNCdEt22BT5In
VQX2IVD2i3WTo2S/uodm6wSe3IjdIPfOQJALcoFTqVaOlQnx+9rQvR5qaRNsF/Q0
08KelRuyPPJ3tI7p7v9ILPEcQ7puR95nro1Pxva324UA0u08YTfRbpIMWSjdEpyW
aGsi6FUH4lv5MQIYjusRF6H5i1fFojLSYm1kcvXl15tFenGHst8vz1MCHVJSFS6o
ioA0uTM1EaJfiOHwNZ4tKfh+PV2RCTbHBN/4GFtaMFgoOJXBaVHL7VMns1mZHl6i
pCqs9+dMuaCvC28lvjFI0nnnetnT60dwWn31Scf4t1ldzdk3aBcbsRBQ1SvAof0p
6P33kwWZZa4OF4JU2U2u7QieEvioL29DbITnesBwP+IRpaC8cJisIMFRwsuiOqsF
87YYxuSKIj6D8y7THAHWIOFDNLNaJUzBbCwvrIqln+mNGKnFceYOyrIWqDMhXXzF
/pGQIT/0co54xr1jxMDqy6GtEtSUFh1YoIcjPB1dHjjcfFu9dhHSfjTsfoCS5ED0
YIbNo3dHAck0OI3mVjwRSx2xRY3icdUSNapFrwx56VBHYGpO2B4ZGtEOrLbLtCnL
1dyNeu+k1nc/1UT0GqXlU0s0pYLTggMeXahDKMc7IUmN1KZdKAyntMcHWUCUKxbd
I51tEZpL4/2Z7FUY3mvOFxE49sJzBLJ9gJp6RX1fi7+0lG2G36+nPh0TC1EuKNW2
xaCgZ/kJF0RuxjCTf0sCOM1HqP/hxn32LWWOGbeITyYVmgxSqGtCb02U1opYwqXH
ftAyKRNnO6JJjCjFEQNfUsvsJtwpwudxupKHstqh6hNwwefT7EDI7KoJfFjyKCHD
8RnVGJBDV6bwGWyN5tirdLzhFVGOAKsBoQABOM0its+9CZrdTEkVUcsAIecvdd35
lZ/ipKzOVwIFiqYayWX2wMZSeVp2eBLHeRfT3VETFhgsGas5nlzJNKD1s4HTwDp4
c1EduNhVqqi2ye3229iwJAYkGKiQ+boeERhMSVwKYA7W0AX3b+Zo0m4fXrqr/GUv
TWP8N9dEfRkDZifaXY6TX34WDskZF+vw32BOW1boiJkwyPaxh0ZRxy7Pz4Dzhwaq
4ULBEfErHtFMxT9am/J4z26Z+ejagObpb4dtkyp4+d9EgI8QENXM+Ju03+OZ7/0T
oo6KA6RLZq5q1Gk04EFi7nAbcdEQFe96tCWTXeGSseuBh43mOAWugEiOPWk8LPcN
GhBvE+VP8md/CwOaOhde3eNr3mtmBiwIjjMV49cVDBrzOzpUd7IGCVFnOsuOvNvD
36XLpK5bKo8SZ+1ZXA0HmcYUCGBaOZh/4c+jbBBGadiur0mpcKmgQ6rdrLiXGx/C
TfMttzoj/FqtmhHlUlC5eYTfQ6BoYPcYsFzScVTTBLFQ84jAU3cbLc6ovxsYAR58
Nha4xkQRYm6+KtEPJPWfRxo+d5MHfhDYwpd7qZCN0XDmwPIKREN4QNUO9L99IA3c
CeFnK7HU/yiWXqqM/2KSD141bjSmajtshIUZaZ9xTPYevHXHnuK7Zdlg4oHu86Qj
RsrUFvsuPc+i5gY6Z1SXcwT66jR1kJLKNtBMFtAs0zEp1M+KJKOK199cP6k+Z1W6
7kIoaeoYMF6ykb39PTKX0Edv0AjNuvXISP9MGJkDABKovVLzt9CnQSWjhZeYm5sh
Di9Ty7QB9JLBqVsGuXQULLxp4MMV4Wb5vAVwJpMMJC5PLf9sWJ/KoI6Z4rv/+1Gs
Wn+ZYVf2de0euA5Q36mW1DSh9Vs/PgwCtHBz2dLeyeM0P4SjbVAClKVTv8MSCRl3
yMCrnvnE7iMIrC+sLGaYcAKSghgO+Q45DcyIN5EZJirwL9pBvcTBhuvcRtdV8Emb
VVC5v2r8AglU4XxtkHj6eefvt5jzMI6WVkNgFVw9g3prn4u1Va1gI0Ou6UbqTFON
SWImOHXPyOvdzKbIz6cAUnJwZGYSgzn+k8DZ+3rXjGQe1KDirHqS370oOmQrpyLk
Qv6ZJu6+wY12WiBIWN7yfoBCqlS8xrkECyXbIL9X9kslZmdMQZSIVAZWpy+alSxB
mdUz0Stegm0ssE4VOWRcO1Wz7UeCaqR5hBt3pQimC/7OoDi8krNFoiBOpmL1CMCV
qJVd5t4sIczEqmG2fhmDcb8KoWCX102WQ8r4G4rjrB+zR7pqueH6F9s+oNDCspXa
TKlkjVDt9ceUoBVKDRAbEfirXlCShpjBYwMrLDpaesGr4yPVQqP57qqYk/c+CCWl
UhqlPyBT1HIl2f5kUQ3kbTZiVwdhXlgBkqADp8mrklETTK5vum8qYHyeUkIvOA/r
s1h2RSx5uJsBO0X31xqK4aaOXRrxPnXqqikMEuVHqAjuD9AfubQNSx+k9Q+k9lCr
91FG6JfevyVRVcme9cCaR43XTBUYvulD51Ho4jCfJDlmByJLVDzHhdNbtr3Lb4iI
kVkkj/OTm07D7fXnxq21HB1AEfjlk0khBw8KifqsNa4kNUsUYM9NiYzShnnrbp6G
qb+TStV11oIWqGwKtUwDPr0pulkVNX2ZzGUVEN0EwFNNm0Vwthd2NBGm55QKyGG4
oy2ejwz9scmhhrVDPZUGQmjmG/wx1pQns8mLrJM+RcY+6iYb9d6F56HfDBM5jNSi
dg441ZhVlHz4wsGKFwcWZ3suq6wMPhgqzUUbzF3ikyaiKemdA5HiVBmZygf8Wpy3
lQJ8RbAgnmfqmf2iRNZfqY+UOlPrNDeJwnmJPgzeiZcMF27xXijFVsjqOu4Cjbqp
Mmg8kAXi+I2vDUjJH8IZqSjwouqHxYV0o9yUNl2DsB+lQCVSHUp7Ojb4jBRRsOhb
n9J3RixQjrdZC/gEpv1vu48DCOZBj7XEssdiz/nfJ6XSvIbD6hAE/czc+j4nn3fI
VG8W4Iimb3XlD7UceAAHGeGY22uWAut6o0x53jg5FeNy3CtSorSUf9YUcipui6E4
M8kMT93/PvNNc6Wo8ERub/VoJEAz6qWGfAk+aCrfwaD9D4E81uLrRVnWBEHiTLkF
in3di9O3V5A7BchqDBf7rQq7Ctmh9pQiQhymCEfgSKgx6YSm+y6fOVt11sMvVTNd
ow4biqedLyQTzmsgeBA5ECKiq1B/i/HTsq0eWeUKANADQ4scsYkErzMHqACmDacY
/rQFf8QqRO8f5cVFXCvSLv/GWzYdS5TDfY4wpMQ3ApPveGbxvuaieDLztWt8TQ+P
LFwzPx1Dxp7i4H3AsxEWx4/uCvvuJUU2H7PpDD835vhHfjWdlJtGxEbjjgvApXhT
ELW3k/IZOpfkIJ+LI2EAy7O9KpBjakcYjkD0VvatHU1C43oaO5yVDDExOZ1E5ZSQ
/B6JnYG09amAQtoWeq5pIGu/s8MpChA00R0eBKGP3cqRI7wGdM0csnCmZahl+eMz
sRpJ/UEQnX+2KJZadpZzBSGCberXu7j4UyLywFGDQf21l5gKQxHlKh0YPMwo+G+Z
wPQwyuAEnVIvdw5+KnUJTz5MtYv7CmPTX308JNjz6HicJbkIGdfn24U50Kef8jHI
cqdgEj8/AnoxrOYpjapLyvcbZOWGURLIpdZyV/jmy87F0/kpGzEddx4VZVAl1E18
FLWfkIUSfvr8jpBAw3j5evW0wgOkmvAFiXCk2ffe5ahNOMlJWi31dBG9ZfBg5rNp
Aas5G/6LL3GqOPLXUlAMBpoTChOfPF+RmeBFEYuLZvaIbEcY0zKool2t5NKbCKl4
HHDCUwpDTXO1tT60PWqoTVM7HNe/zehMjYjFF3qI00q5Fb8iXi0ajwok9iPle3q4
TzDqXt3cn36cfEyQGMhYrk9WidWx/Xvqbxdl9YoYA7vfG9kkMJF7WBxJlJJbEdOp
4F6YxJrFamtgvsdeAPNOxidqthFB3Rb+5tAiyT6zbYpFHHvay7k2Rr7f83u/0ZrJ
SGh0WGSv052L/jGPW8DUxX1xEX4G0UTO6nXYLeRYV0UvScTMTLrTcRlcM6lIS796
jGV3qYucD+/GFv5Ex+BTwrEzEVIFQouovuFQUzgUSvFRWsGEo+FZUajMoBYiUxui
YaxiNx/1WAKKOx1de9X4/akrXy2W3E//b21SHjcYu65znKFuG4Q9Y+M5GX8WBdP1
zVVxd4lghWpj1zsRqmbvixl8UVoZvJEBbcfU9aAbRnAty08/g0RCjfEDrm5rPZDf
JUkeLP21bv+dhW+DoYFBeFU3329IjCnHTHMa3pcrMPwicXHn06i8cociOHkvk8GP
1NQYfiT0RbhXeSk7yu+uISchvGuEKB3YXqLEOZ86AyogAIgebwFH1XEd91njjbLj
Ce9S0bM1fxgCoHIadjYLDyuXyp2JYswuHw9H80UFBQPl7PYCwIuO885jw35UGh4x
xRbWS474vc00ke35l0Kyy6EG0KXdbwM7MQaLwbh7lskr0t5cLtJHxhpee3sY7mko
DHPcMGsl8AMTWRHhlMcX7YOhPhwlYIvHmsXMYVOcXakExAoBuNCGyOFS834XOxrC
JVwNECJJYQGSIt95PavbTzq2++wvbsDkMz0xVUkSL2iZhUepDV6ufMDb/+88TX7S
K439IZTSqw8x5PNWTjVU6pkfgqwu1xgohn4QklPWL7kwWslRg8Houc5cddN70IXx
1n+vevsFM8wttucYISd9VhTguqiEaanzXBOZmKpLAMPicY6qE+sIHf48bE4HiLs6
OD3SqQ2kPjx04r3/crKFz8EPrzwmrjfP/WUK+eqWGtR6Mzp1cchl2zPKPmw2qYrW
DNRc0YeiipFhQX39QGOJ4bpGW0Q18gugQVu6I3Nex01KH+mO9E1tXsuP7DAScRtx
+VNT54TIXOoCM4AbgeJz7YKKrtY5u/TWzZ9r4t6BbF1yAI5T89Hrj/MIKm4Uh3cc
ngLfX+wXn1kH23qECT0InBHq4E6iW49LcrfyIs34FVCRimwm9uRF2EutwD4mFTCY
LKosBOYbuqlFLJ+zvZ0hyJ4/uTPtvDX/5PxVwluhSPg20e0nXtAUBs3NNhPCSFXj
b3Za++IXBHwFbyIK1PV5rKS3A6B06d3G8qp40ilwUVNnZ0647x+M2+q/g6PhCZ+l
4rKujsYmzz8HFKNCfVrgO8cvn+HxHMMMe4e7FlVtJE+rH96U7rcBsJhhuSbDAQEz
yTx0MkokZdl6bmb89Aw1LuiMkHVPXcNOkzqkt+Kl2kYSVBa89beMlNrresZ8PdkR
2X6UfC01dDYf55FO45K5sydJ4/Q+dhEQEWpLTo2tivyTlVzkUciNFrlJxFgxB019
GnXgIjHYDNhh3kmFb4V1FhYOGzjUgi/f15WnKUh0Wzi2UaswHKsMVaJBuShN6tRT
S3vfEl0m7qwozvRUWBY8hZYxv0FGuxeLunlwoguHBuW+5BYh3+mlBiYkCiPFNHw5
w6D2XZ/WvTYH+akLi6vKorNlZfc41MM6JMecly9lHTn+JoFGP6fSjir3JyJ9WbUb
UWgKA6pgqWaYwuAwonKLxLQZuR3B4I0aAIjsu4eHayIkycX0McuQBMb4YWAgYQRc
D4Pk6H782AoswhXhK2NtLi+ANOI4wT8waNvhdIFnldKRK+NQXQRDLUNkZxjI26Ps
7Gxm/UwpXUbLmcfjUDERLVIwNEUKhU4aZ4+8Zh1QBk56Einus+pqSiBA/oRSdZRI
363TOzaohs5WHCvEWYmnMacd1Z1uqSYeIG78VtMJKw71t01Yh7j1qc7u0YCyU49c
/THxXQzDkk5i5UrTiGNXO2wC8BBKZ1+Q6FZCBPGtsyfXMH6VDBfhgYCrS/85YKdR
iWPBqf3xfqnadYeFcYprP1dOjpEVZMRTC5EDxUBbEaoonJOAc1qtfbr2dtrmgZyp
rgzBuwQ4PDMmSidfncA/3qy7QV6imZHpJBg8C+sV8e4PyAlAZM621kpv52gF8IJe
6EfstWLIsjWN5Snm/WLhJrsWGsEFvMUL6IBzA9cN/pD5lyeOyG3xk/VDkViFLfen
QtA8uAuKst/0UIOsZs2BZVIUUGTO/gGScBvPI69Ni3MXA356wbKU1IZy1z2kjX5P
U2TvmtcOKDdFdDOSCOja2kJHYZjDBs1+EgGxKXOSrtXqceMER7I1HaxkPpHvcu4+
1kuZ0/NtdzQurINvwS8eWUMc4smvUJguzUcbqqoVDZSnOtyr1vS9xVmmDyN+8TMS
698vrlrDw0h8X2jXF0DseCrYBRNt0jpHXowXWqmKQOFDWuwIbbxibhvD/vYNl0MR
YRTTdrO7PndPVjYBHOJp/iEwQPFgLWyTQZwAQiWDKq8KAuux+MJBv40U/qJ3cTkl
aDcUvUI3tcAgf7LA45PWC07AQVZwsn8z/iYiWbw3h2nrkg1ZjDIFVweMbE69SGAC
2nk1qiLrUu7GQGni4Lv1pqGNH42A6STYxf4HI0DXWgPbiCNjlcYc+a/SmGXeItte
0b4ljgEklJVox8hw6XqSDUzzWFrYHkQ6EPbUFErksL+BFy3vxU3uv/oVfkCLzHoB
R5N1hQtcTAYqUbXTMjquU8KyVHL/0i0bq7pU0TUbEjd0ThjNlbOt0oh+fgbJIt+8
mQYbxei+O1yIn0sNRh0XQxwxHtrBwiJ2AFFhR5rRE01C1bLjzjLs8jHZ5cdfN8G7
5D73GlKrfUb8WiiUVyazLkS1Sm+BoiU9VsYzdcpNKYS8c0V7adfffNWVIBnenfUc
Ffh3nIKp4ZLoZhUgFN4atJgFsPqLifRIm+223ZpHUiqutTIEwHPcpRbVrrBLLPJ4
T2OKqZcLcGeDkbfqO8QyII8/G9EBb1oTq/SZsIoWzYEEhU0I/JDFQ918jWUJT6ER
5Dvti5POHjieEqQCB+iApyk6EXjEAxADCLIu7E4Gjmxskh+zClEf5rMho8++20KI
DkRqRUdP0U6/BWF2N2LhxeJvJpVJQOGYNcWgxyjEN70Gyc+0n8nV9wt9ZKW/JsI0
U0CGV7m0uoGby0/Hb6BIkyJjVVIDxfukllpI9hMlX3/2f49sBpAsmQ/eJvSmioPo
yn5g1WMGZMBZ6wAgrgZ7MJri7FomLyjD23aKXUnbT9MzqN5ByoZ5lNtvX7vNjJ3f
XqL51gAVKW/Gyb/M7WEz11mRWjMzHN7oaaOxhndII8Y0nP6dXe9GzfiXMBcLNvkd
U28Jvb4TDRRiPRwx1NoBdvezeT7eL9PtJwPY8T85bmyx832C9l9EZXdpU1sH4rJz
RcwdRgZR1SoX9GXEBdSAaK6TggrW82cLzF03dpXqjCVQmJTvMeNmm4oEdtBc1486
Nw100JvUF8nKYYC5W9xtg/Q1nZvFnR2LIpi4pHZkUoORGDan1D+uQijMPcKj7kpP
4YytuN9qLg54p/dW5NJP506/CuZtY4khK8b2ZCRBxgTjrg/fWFxgTJne5IL6DV6a
RLGwP31DI1bDyM8Symcvk2gRYZNEXzVS3Dq7wlxbtHALtU6K9pzEWnf4Nqz8o0+c
h5rjGk3ax+RWajDgVOO7HXQ34wtp/16UYgAeY5p5WVAWDfaRl02jRcqEFP9sTShp
CuzUT1WW1KXrqrCU9JJvwtQFg0KfJeVS7h7qN9jmTvG126J7IeUEUL7rjSgh+sFW
N23l7NDln4R4mv2i39gczhGP8QfS+Ami19mwGsnehzWUlM6g8Ajga2+FUtCcYxE5
BCAfHBx98Ow5MwiBQybbX4hSGO4qoxmnF76mVgX9pUSf52NBA7HlY3LpRWe6yDCQ
XEXi6yiYqwpC5DUBcSf+rVaMVT9UMfZhhj8ymI9EKNrNDoE4eW9TF+zK6dZ6okh+
rLIwKFIC+Rr9x3x00fZMI6vzdqy0tgGNySLPREoGpDD2qMm3wq/lZbgdmrFuV3XV
d1eR/1i1O+b+KfCWWUePcEo2DKzLfdyr3zXX2CRiOSSpHN+0boiNYFyQeaXO1NL9
WExYmSPxRDWtwJhGAdbIqJ3PlTYpAsjTBZ7onxiXZ/cyFWPcO7HQ/3o40QItQznN
AHs+QMhc/PegllMi8a+PNvFIa0nLO8NHDiPvHxwG/HHfM8W2+B+fipYeZV3kV5QX
4y/PbeM5PDdOU33H6Rl2zRPSNQTQtuv2bEk1O4o6CRNaFL+wlW5wTlcP+luFezEA
40yxuevletjtFgsmCI757TtzhhJMje8Et5ERDgTy3yA7fDJc01YQafk5yIsUHhBd
e27LwgI4kWOIyagObyDfzZdlntAkHNtlY1R0cXTF/SO++zVAyV3QGzcZS3woIlll
OHp30WI0Uu2tcp3VKHVESD2hn58RVbZ4XTGwEr1knNZSBeialj6xaSQfpfgw09Xv
18/ucHVcPL2Zh0Jw8WEx49Lg/cUju2qiZG7h4c5XbXB84QCJn3euyLHPVO2L/KBL
xJh7x/xtBiWNq52OEw5hzleziOSx8ETB8OcSQeCke+KQDip7vvTGT4r/RJXv3v48
hJb1b38pWo3Fw1lQij4poh/qe1a072T6wKQNfgKvaNKG+mOFAmT+rht1qZCR3rmK
CJCvizpdz2FAQKDvijOFB1KvIyF8cqpOMnvWf+d9pTd/96mxGZGDxI8isZdVgKi9
nv+q5pjrFsDTsBDCwVooFNWi7FTSVF67UFVyoKg2Til4nylbSMwfJv/NwhCgkW/H
q4moI7guN0Q5u0+UnO53hxgFg2gRp8sIa7YckLLhvrd5SghSlbb1N/M84ehP6oWP
X9w0BHCLlbWRel5ZiWfWFd0vodeEdkGBmIxtM9TAlIf7q98wxBv0FVAE+eZ5Px0f
J5rK+zOTpztDH8NmnQ3LZKkxBb3bWH9rK2+9iam8mS5aWG7rEHnIlhJYN9aZ+ldd
AA9PD6rgJmE5PG0xDv90AFMNED4BjqhXW44yyf/k/FBd3ZHMG3/9TIsRA3EmkqtA
JUwb6bEK6tkq3ezSWHhzhI/O3AxLBF/XGbl/f5RdE1jZpx8ik/YeeI2b+M1bt2vD
UF5t6TU/fwBPp7BY2t2HUQdqpgL7ooNvV/CuMOghqqZIGe2UMdLVb2DxDp1W6Zt9
W7ne98MqUcWunGgFMZ0Q/ghLNcwkwiV/j3YFBqfFsM5GGVRgB7frzijXDjBcG8Ar
Edw3/PM1J6+Ca554VQLBgHK1ARNnNv8CUtXd8Zf0OaZtkOallOkzFbOSXCVmnCvo
PzQE8+ORM1UG9aNHn5athiaDxzY9Bs0sCaV4F32Pt9PXmXWSeX7rhhB4rvDJZ0uy
lnKss4c+/Zm+Sb3POcP45laYGYIIqRMJ5uetp2WFxbkutJ83Sfd1yNNaQ21D8OoN
JuXHWvORNON35dPbcLS6LgBXMpXJMIDfhZPLm25/Y9AE4eH50XaOOK81iHZntLBV
toKvYDJgiYshOLqYdOns5qYGqFGdMxByDb5N4EOA1Rz4l0vt4CxEH5EBT7/cbblM
oRUnShY+a8OFG3ilzDQXAOBrjNFJOErmc3BsNVNBH6hv5Ym9aedvRUrJzGvLFWxr
HA/OFTuZF7zlZI+3THaGIiE+WNyxVRsYKZZqdjT3zt+0xxOmDOIEgMwvupdUIdEC
R+QMu1SlWmv6JndHnyITy+Q3IA9kkLbBE8FjbNFoxCNkviswppvIZgyymlLIZDy0
8DDrieoGeWo5J1U7KFEDHB1qggjYoRmUbnfgIf+guw4ReOWjgloC1i+p56YD8Xxc
Is3aIYUr0iKISLb883H/VV7CUmodNyHTNE3qKfRrI1zCDuG6Vv3KEPAd0BhLOrAS
cZy8LgdnCOTGcqHVUt2B2zt6e0ar8KvVmpeefZ5/1neDGR7HaKxdLKys0SBUdIiK
Mrj2LPJzUmzTFFhKu/X8WFIgKbotJ65eDN+0O7YD1a31q12W1CvFmafxLX01t9Q9
vCTiOOIbVFmd2nZbp9HHEFlnfeHczM/JN8fl4UMIQp+hNFtj/n62UU1xjnY19BdF
DJlobA6gek506/bui4v5OGQ5LBJm7ko1jOE+WqG9JopOXJwmQN9pW+oVZ52/UrAe
BrUxaHGIIAV0oqCFspwnc2PStYhDJHn5uMcg0c3fidq3kBHRCzkmzcAHAm7wni6s
UlOF0b9MOxZCqbvmnz6RfiulauhKNzo7gEuHVxE7zPwJlesegzo9VLRNF77I/uh/
pCQ8aGq/6BlWjSzH914IB9pyHrHdRSe5r1TUV/hMB019p21/n8SoYDWb+sqeiBws
Bo5bOd42woB8A850RT0ySZjVRxFvND4vKS+GrOk0YkbBy7fUkBCrqa0UU739QR6f
kohmPStOUklPzAeOxg47lZYzgjiFnZxv18Z810YCIR+epDYYf4yrtUNsO2DguqHP
wna4zCVMEBDIVS1mIjlCPpGYf61H1WLOeGOO0qarYg0GV6l/33qKFNBWjgmyO0/j
GtKeUaB7xZ9Z/s6oduAjzWUE/fdi5arTF8lPtGhoZmTk9ROb7qkkDhTxS+YmrmwP
e5ycf8kFPnIIERM7v3hMXDf7X9+S6v93CklUQj2AEdgQXxtS4ey1jpSon/VSqxYH
ddj+DykJW+LvTX2ZoOenL7UvxwdQcPH9UXvrZOvvPMA3wNBYBPUybuioP4599OKn
iVWi1oBbRKd3MpI5WL55QtseJ5n+cPzVU4VvxRMsoOUbF0m+OUSlThCnl9DSaNEI
xRcLgXFJ/v6ITqDpMoY4FCPVxhsy4md9FxvzV0hLm362lJUeMv4ORAgYzYsc1eOZ
tkSjgmKiTW5q9cX6pk/56xssySrS8UTNxis/e8BG7AlfwFa29seiBU0t281mVtZF
f2YLJll593gi6EMXB4E5Ou/GDwLX9muUGXONv/opqwbnZ6impH1X7Tss6OYNXlS1
pw6AaqW/68wu7z+xWVnis88VLJHGL4VJe9cWclex/WdgqkH72+gMPKVlU9QE+6Jj
gEAXHnakEFexjD8It3XFB4yt9kbQ1f0anhEBpy+Kjtssv9IaTyMoYugkcdus7V6c
IG3tWoBMVEsHOyH1ewL7V9S8vD+MryU+iVlhz+LiZ3WKZayv++pEdbNwU4f9Wtwq
0rQTDYT+slh8zDhPi7j48LKVMpNZUFdkw+/6HM1M4ninzws4z6NNhmt6lpo0jSJX
gmcTZQ4OLiaguhATY7R0ymBtkJIYnsmoL+IQOvrb7lyEJiQ/51GaWs8Amiy9Q7hI
MkypmcHLGNzPboT40Qhlu+iCGol7qCWvx3j3fMfupBtaOI3Pynns6ujjlOx3UMxP
fKTpF7gPMKTWbfpNSw4A9mKV52flFSBsjZhvGMH2lVjkOsshub8xPupaIz57v2xa
ZEypBI61oculUfadFEfouCMQXIltZZXPXpr/er5TSQ0hNsZXSU4gNZq4odo2vy3o
bDbeQQgRkFsj1KRFluLFin4WzgZHBtlkrMTmV2uSJVU71/aCnMeB0vSQ/nNo0xvl
A2zb82p2T4bvK39jKjMh0b6MmcD7cPJtmyalzGI2HO3+5ADp9wWrlV6wCtzBSo0r
RlCNlOIikN/k9Y+WGibgCBMnHJ9MK85/g+9L0y7ovRVxlVH+hTksWFJmddAmilb7
icpTlPu+8LJbO0jYEpMyuAZT3e3zos1aOkpb6lNXcKygtJiRVx+ihBnpZXjNxZiH
5BcjpjXlhmBhFuas+/S8zCUGI3BoS5uEQNfBhl9ZS36vBIi0Jjo0LCjLZfwqo2iO
tWSoOkv7V7EPBWXBbtnwNz0WARj4p/ZH7NOPc5RbYGU4jdLefamOUQcy5ikg7cAy
tSGbKhWUG2U2c+J73MgJa4BIUYZA4tTvWbkBOUKgDI5qXATxiXmAJyza7C4fP0jW
i7ZPJHlkPOxOKaVvsLaHCHjPCJAq1yMmWgR3h4MA6NeVCr4MSNKbSEsmw4r18yIR
vdxo1+BhtN5L94q77+vLJ+PmI2L/qMlki7rDsGj4gykFvtg/SKIKFjsFJYHZJ1Pl
qwcRtnyvEeDLFK4hZU5FakOxj1TN6pEOeADynUpZ2O2t+XHRAoxsMswAcLLTB/vV
owqdDCbWvo/uY69/+GTK+/wyPB/W9pWsF6WTIO1XJmspA25FhOIH2ASb50Amrhnm
cy2j/HS+n9oWdKOzznvNq/AXnqt551RvJk5oambpzTKJ9qo+pw+sUCqkE0rOMS3T
PdBdrMhVmTGFxpvdR5CSmzsxg4knz2hiNEDmjwZuVk1Zvg9H3Fht/4n6HwMHCwRN
j70pWrkhPkxbgttVYDNYOkUbMATRMFzViANGgVvpsagw9GM+9WQLxHmsjuP6bSwN
eLD+r1sAssy/m/yumbHoME8vQQpnHPcDFG+bSFdRn8snLAtYHHBPwbuJSsNDMJtc
wVZEpkukbOjAD39fExlKruqDSLeRKgiUSFovEwu9nidRLeEhn7l2AxnccxZYZEL/
Iw7w8vm5IUb3QUlhSPqUgjMWdiHaJA4yDK3Hi7k+55x5044I+7L1AXK5xkLOggnb
NZ9ChjpP9XUFafDGdkfoXXJ74iBMSVOK/YT123lG7Q3imkEDCnfeLvunjcUny7Zo
vn/+spQDJ3XjAenPZkF0j0yYpDTN90WFivjj38bQfI2zlx2NrKJ+tfXoyR5FeM0L
RcztZT0h8qbXsune7eTGGPstsyfeSwOCAHlz5ZfN/sXuPx5P9dGgFjjT5CiZADlv
gxqlyNrV9xITip4KGZOEnto8Bz6KFscQdpNCopxoziqGd+N1EasfIs8Vu/rpMVNC
sJviSquOC7ba1JZHpaMHHt+FBHr63MGGSiZe4cRC7VV9eoSa98jnE5l/AS8v6021
5ozsLKJ/mp5q8itvvJ4Z4Df5rGBP5XYmb6YiI1wqrQX++YX5yZ+mQkMTy/HHNbRg
lH3q7cGlBU6d7cjQ5zvqlJHLYN/JMOEadzDHdPb6CaoRsmItG4JYHwBv1DEYMhNj
rLq2qw67arx6s81N6EsTQs33MxvDHpQFbhZD/XCgeGSfp608MQKGVsMLCRl8FQ7Y
KWTTB19+7DMQNB9PSxaCk8OspUekaq4A1OAUuXkO0LzJCYEnPPBGQZlYhmOGqbS4
YVbSfYjscQsh+jM2wukAC7DbaljSrvkjVBQ5wpUJvqx0IBol4jjo3d2wX1iOQiDn
mD0QIH2bvPtSBdEI+DMNMDc0Y8OfqDROnOGY8FZshy7h87GiAyglSZ/tAKewz3N7
Iebk/siUVE++P1Th59my021n+PjLrRP5faw9X/DLgTQZDFvrDqSPPKE2Syq5Wnvg
eJViZX4weTawfet5Ot9u3l+JduW0sRAVZ311kxyRmCYbZU0ijkIEP1CSJQccqGmS
nSZYzMvcUTmjyzM8K8vssgHyFomUD1Ic7nC/F1yxpdOFB0WVidjxyjkeopyh59ZN
q08da1Mv8jc0ViIooS5xc/JExzqQ/9Y9FTF40DkEFUengUe6HuK9riWjSscSshel
+67cZjR1aairMi0dJ9CGoK/+Jo9AEKUvE/A6uxjcYDqHODXVYW59X13L/2t7aoB4
CyBaLm41qhfoXD8lwYNHIJ5cNvrVP8+eq2TIRN+38XvhR+8rEU6KLmwksA1BV7rg
sIPLtlHZ6shoe2p6XVfZN1F8Y+F2D2wwN7nGN/Cx8NZsQ/sTuC8AnLY3sfPC0E8f
WbUiNKXQlsn9C+Tvx5nw3yXehessgD04cE5c7DQrS2H+BJIulhmp5SylanK4hkYG
0/bYWjxTxBqF1x7UjYJBZQnX4TUprx6GebEYe4EWDhTWvH3jksUMJgiCUw0w0wM5
28WzxHpbtDzt523h0L9EQtPK8nXtJHrQfYBUmAYJgHydYnf0+3wWCxBAYn8aPqQz
MmJZdHbteDya8u0tHyiuA6oqmOTiJG/I3qQuwo+WbBGb8TR3bsi5gfMC9XmKdR7n
4Rp0Dsms5scMlVEL/OIIuJGMuprwi+jYG/wpcO2ZU/X5vQkNjHuXWcdJ7ID0vVrF
qjzb8IP83dPkgujsC16Vk7g0BwKaMqqH01/aLXvvEk0vr8BXyL2+1a5sgMnuhywL
pEcDez/EsbERUvl2REX3YzpdsfaaFfQ8ATdb4JHkY8rJst8NJZUQvA9VruqyQXtF
ktOx1c9gTuJezBN56KZYDBQkIIGb/vRCSm0DsYVe9sldyqdCbjhNkJP269xuYwqp
DOf5w8+XEheMRvgz8hWzPn11FXsEstwKM+nA0g4mUUnSBMfRceG0SaPZg4hZhF5m
7HZQNNUgD/jex2ml5h3Y+uk+29jursvdXZETThg3fRm6AnIluJvJtV1y5pAwagkJ
jIs9KAxo1CvlO7zWmePI/zEhJK8A23xAUo/G0Jc8HFkGpdIbJktFYGqvefNQkxay
2EeM6CCB675R9VywNZI56UOooGljG0stf5JI2nJh8MYrw5TvgvlcHvd3YTOXMU3p
VisbuuwvgzCGzfLTmjuw2m0qiYMLY2MjElVO5a93Wevp2UaZ0xcsCCW2Z8Lj7sA+
A43afUf/2e6e9RwS0DYdRQLO7oBKnaxMztikRliv1tTXgP9x/2ACPUeV9Rlef+3H
vEaUoEl9sw6EqIhkQboD79hiMQKtFLBjfIsmPTgsDUaGX4wSJgUt9gI7Di2AbsKd
G/lCgHrAWP4tlHpgzX0GaQJ/tqXiP4W8jVJeVzVlfbMuQ4vNEFJWYZ7FaY4O86Qw
n62iQGoQsQKND8sGrbdhQpoA1S9H0VFt1fm/BCqGKLz6uBvA/fKPRVG4BDrhnf1k
FuBiJ2xihH92MFgZqTQMzAs1fjXovl2U07NT+DR+CxAVdiO1HZZeBgkiQvaV9ab8
tR7IXmWsbaSp+WtVvx0t3Y5DA9KzsVU8dV/VRqATKEGnBZ+t6W1DL8lNUIEZcaEU
EpsRWIJDBishAZaTs7dkGlJ3GEQFr1n47zVIDxl0Dvvsro2+1Op5InDsJ24yGYvd
bp6zUg7tCZ68LAq/7tB8s1bhkl5EtJQqaF+UzBBXENI0ZGtkvcDjTFkiWLdtyn/+
o7+tskIWh94WGOP1A62fE34ylUfnm+M7r/X0u4Xirq7tKB5tHWebzTPdvDZjhiXo
8+zbOaP+FgXxUY1Cxud5G1Fd8DFwcCHaqC1j7NuD/MAiJ38/5o1goyDKfa3cAfQp
gF+z9nSx+bKxkIeWL6/vamtnQsO2nNdCsUxSIFBcz8r6lXjte3zGPKAXE037FFmk
0yFVd1DGil7CW4/AQSnDoEUWRvawMwEYWZaFDBo92bKGaEIy5vyj82GN+43plItd
9a4vZtDvekySxuhmHtvrTWE7VLuz+zcthRisF/CF68ettJFv5GJq/hVV9HW/rqQM
57aWjjR+Gxp1iuyaboT0tZ3MqyZi5TQizlBjcaGbQ9a+jKdmDEiJsEtrcrBAbrma
3PZeuDISbneKq8y28F4QHVGPrNJcwQ/tABiI5pcJKRoYXJfa5PJxtMsXcXDHQTh9
ZnTTSnPJoRATkDVoC76A60Og3+Q6yiKehpzjKRTVelwCIb1HpH3/xFWwhjfE/P3b
KAzweW1RKNIqPwKUiRiDMQxK6A1maXiSO/SVaXnnIdSFb2Sr9q9iXj5SBsOWyWvv
ZqCaYi6dfJNlRkZhhi2RF5Fv8DdY6oQ2abiEha8CGV5PQN2rrZzuHHmA2yj59MUe
kfLdJKrda4I92+uSFxGLDSYCSNiyE2eJlslmvldxbfX9NWDnQ6PnEM/17kbKl560
4tVhzT81f/n2i8NW8Gl+lVxTfHjDXbcbA6Q+IFN7cc56NiV3ioohAeCu3E/wLzvU
TBqpfNVowgKmMJjJqKe+5IcXwT+ztEOqzndWUkvU0czcu531dRGHbJ6DnvQO+Og2
ousqjXUItjrkHcYa+gvGQalTztC87g1u7Xq4Z1TrS2u40RhTEKhAzg/zHwjcZq75
iiWwqH34LL6HPAhg5d1kwKoeCvP42e3VttPFxkCv3mlPdMyMkFEnNtkdr5qFrHHi
jb2DGZay5zlm2lzZDOpidPkuc6N3pgyDTxkgYeoJXuMc9r7EIIzFrHM27DyVTbSk
qxI0mNa/3G41WD9GUvRvSMWT9w2F4PZ0jYz7kcmtMccrj0R7b/irj+ECWGJQ2mqj
QEBcZSBUUtjy8uNn5dtYj/LJBL9fY3C6VndHc6ReGYjZXzp21AbLnNh3/GWqFA9W
/4wk3auraP9l4ZnKSkuVsaNkC54fXGdMMqC53+QIqF+tDiGizEBeRkigo9ptPQym
ckCE6fgjZ5khinUG8c6Z/nU9a8m1aIv7RuztnNDvR6lUmX2ezTsG75ug/q6JVw+X
ePP6K2scnK8wPe1szwhbRjoSyJSwTFRu0ml/enRhUKyPteSP2GQYoT6C8bZoAbzJ
ADkos8UNzVkietXlb5fBG2/9G/MXiSJAf6rSauFnBppAdWGZ1iDpRuFMpQ+yFMlw
Zrx4Y03B1OFbOMrr2MwUEc3br6LMV2cOufGamIB32lARPEmKY4npEw5Fh9n3ajsd
GXBKiCxdjyXr9j0yX/i6WF51hKNTRtfZpBl0oYitUk2guxluCFG/LaZw1x6F43X2
P7lPZvKqK0hMFyQCag4FmyQdJLl5i3/njnhKzvOHrpbSUbDC94sjWrmlncHlcQHH
p/89T6j51TMKkIzCmNjn2SbZkgKTKIo9CCwARVNB52ygJtHR+YOOd31WLO3SEbEU
w/JPAryA/Cws060u4vE37BOTtc0sZhuFDPDpT6NOLPlwSm6ZD8y6SROWRWO0hGiy
ItVZ6taQhuXLldjb9ZV9k9yyc6zTXqyoBv/tKrWlCcB5XUPmL4QvrDM4P3SHzoyB
U83o6iz/ET5twjXEM3ilP4jMknxxf3XrI2EQNNfX4goHx76poozIlKlLi0EFgK8K
TRTSdOr8VSIfD8pM0p4+AkfQnprlpJOAnoXjsevx7XTfJ+2cy4++QAe8NZIozWUV
0LL2uTmDFOhon0MgZxjb0R4qMCc+WgUcRzGenZyE8z7wtLD9uFExXnGNb88gSd4e
o0UsmhT90UgR18jxlBdSGH3cfkCU8TAzr2P5sH6Ozhg0gah8Xob29yB7kn7k2Xur
ABF5wHprMzxRD1mDzJ41E9B/6mtxRuElGgpfZH5LejVLWuE1x3gyxalSY6treY1l
ZZHnS8HCLg5Okyqu1X2VUB5SyekNFJ0zcS3kKwyIU0o6S6w1SBy6BUH7bvRV+Yf6
aFEN+baw4mHEremfOX+Zr3aIkHPDmM4ge6+2LIv68Ckua0+i+VDSSQARaxYJ0uvk
uDKMtc/tPfzvj/aZfAspk+kXBH/I8xwsj2jYMPKGN7JrkZTWvUKUztDgC+eyu+FZ
MaLVcOXk+u1usWu/IvvGu/f7VC5IAcj4TboA+2Mw0lVKoIFIVv1HmB+GRfQB+KFi
NzP4cFOquH4dPtquJjxX+Bvs4hfgUAsX7Rr1yzFRbgpG+q3VsuANJFkMajxPmC5H
ZaPfoCIz+31rlGnG4hGBTr/Sd8ckXpaFAyoA24b2YdkAyErD5Cm3udBq0Kt5w3+O
mEnFYylrrT54AOjBiRJY0VSmf43zchPdq6GCcr0aW4Esuo0SvLF2QFmuwaOJsfVR
iT+bVmNr4nr8gFKTHrfHVSd1vj6FdZ7O03ocIabLSvpUinspbeLItXxwdtBlmG18
rF4UtiLtq92wDlPJEU3YCPpjEthvIOi81m7NH8FRXSde3s77G8SWA7aNDsb24GVB
HIIKIT4q0Nly1pgZskXETXYuUvxzpmom3P/U0bLXMCut0W2J/mLurjzylEb3dwu9
jU9ytbaWmJGkrJFgq54o+1e7vnfA/ikSQBNJhvGUF3L3NSe3luVr2xhXTBWhxoz0
VYvqoQYKRVOZToMsR35hhD28Tuw9Oh7U5vLp4kPh05CRME8MdjgJfM5QObvQrPvE
pWKUa4PvtzkkZmteGRdI9Cl+nK/c5GIfnk/1KL7qTkRF+s9q/2/Pltt0X7u6Wicu
rmiSsufOHRDu4lnLifMYmSCzfO1Qgxt3oWTHorUVRVSXjvbG30JA2Hxn1N9cDEY0
4LAwwiinAPFwgvKZJU+BvoAL6GigXOvXwDQXnf7Rdir2/eKB/2kkfaV3zFlRrnEG
pxs99mhUi07OFgJNDupW68rdWVDUgKTEroq4mPVxs6GzMOgB814ZrhDSHvjR+ehk
GNc/AKedc6s7ncAM8vgEYKwH4zHWbmyqcCJlO32Mie/b+dKw00lVPnee4FWR6jUc
Kh7qaXKAX8UWP5pOshARJ2jVh6980i4oWn06QfCWPuzzMI2SVi901k8MllOe2n0I
XDfFVAKglGJ4NZm9T7FXfOjM6j1GqE8mIYox8b2lPCKJSUFFHEaE+olUo3c0ehDy
6pRoHZC3D8d5+QNybBTcuABoHLU8Akp2r8ijXhRNVMi76CA6a+EzOl3bGyQD2lo2
Urdv0E7NcwVxcpEih2mypj8SkOsy8rl6aZaCiYrKqF6SvKV35xYXGBr/+0G/aoUV
XItBilbXvmEGiTIukK4k3XH2myIVJGLetJpdxVXclZOg9HVHRSWn5vxe0WZoqeN0
x7o/93VhOXhzZq463e28Fj71UCay0nxoU/V8E6SGFUlIiY9Lge44K13NUwntbtLE
OQCcJd74EC5+yzYMKpr7Gy/ZCfYqMfoYU+C7DUltVx/HXOoJDe/sN1807vVWclvE
XflG9nVN+uUQO5rJop1Ms8UcWKfIzNPdn/t+eA2O66cgAiQWPWpfswjBUkTrhPhl
DXF/RNW3VmU4e/C4OUjsLRreu9TQL5aZOn3BUjWGm0fSqIkPliEmGpqLSgtDo2UY
oKZ6t3C3jKPYqRZzd58ttuodu/T2IcNttBaorokMEVxCdaoM8dE0zMW91tIz0H14
w9KHlb4zUxLUlftKy7BNHG0WuHLUjRzAxRVXOSDYi5XNUU2rNTBiMRJg9AHsva8c
QaYlBFoFRNDG0rVqWwvUrBV87LMajxiJXcdqgIkBG/liBPoWE8lEVBRuxv53mNEF
+0ENTy5z38a3VGRKagZNUp2uiN7589Ge9SoUWH8FKaImfw4gBWy2iubNPxmmJ4UI
JPFskW0v+ji12jwi04uUvCEF1tmBmWizs4djhgrxHzFt7sz1Kx1CuF8u+b1+3AP5
DSkiCXqTAv34iGbJnUZI+qsQFbri+1blA+XhY73ES4YohawN2naThebWjSMjtfHS
IoKjfR+56WD+Ls0gP12A9CJOPFWFGQyOdnT50DGwJrpOjvpPW4xzaL9ma/OTkspR
O50zv34ej1w+LPcrzrAq1hIV7soB6P4JhM4/mpyEkW2BfPe3//S9YyFZjv8jiSZB
AYjWN1gqfyit8d9nwL8XLsbj/p4zx0dp3uAMCX6LD1cll8Swlj3XPnGUX6FjVZjV
OIVcY5N8E/q0UTg/ZY8qeI9JH3Pdch65u+A/ev5+4mkoXe9R1v85Zv+YB+x+456j
TJLFbXLweVb8XYj8D8KYd1rVdYgdC3TwpauUOW7sDFVVlT4ZjwJKQotX/u+G750D
JvoY+kePZcT49rN746EI2DLnDXSxI0eizZFdLfulLitldFDsSBqsVMdI67/3fbDI
V8vrxufdSa8qafIGBCYI/6X7wD5eTfQEwcaebcukjLbpiB//xjVDT+2fFh76pTAh
ZNzuz1g+tYDAT7xwcQAh7jQ67sV76Bubmpxqf0iytjXGD+SXG8Kb2mF7a0wlHM5h
C2wdgN1hFDHutpqvATn2TQ/ozKDQSE4Rg7pDDgXNeiK8cotQ+h/Vz5+U/Dr05kkF
A8ETj5gaOdTWlOesY7noc7cJngiqjvYluVGONbgVK20C3UNGrHriTSMWYS3gTLto
I++iyMngeL5YSAC9lkgEcGVKVbyPVrNbkPlvXp3rLNIhQWfmP4Oju4bc2ppucei2
GSe7b28Za4tuW2b1U5ztg+nZ1JUAehOkzpW9fgdHVTxGY4xHE9l+JVUGms1a2LRX
CxMExLVMGZ9HarOlRGOo/ylTxGBKtscetKiiFCVEhP+PFS4XmPATbVCDe9KLLe6u
3TZUduT7FBpYhxkE6fSzmxq/E648UUsIWEl3pQmELnIm9rbpqLEhrYEnNbFbp7BH
FFp/8NR2jjk/91XT1tB56f6FyWLT/yInMN1ljEGm4B+wYUiHoNNvk8e2TWC3AS0r
8N99i75QTlpsiyag4FYPPXsdT3Ocl+g0cH/R0a0q1XSarGL62LUuQIuvLUgG1o2b
rEHNjVJNnuxzBQzg7Ly/r1VIu+ZdGob0uUEOs/iT4YNtxfmr9g2mG0uUn5IyYwYc
l1nAHnDeakU0FnHSqRMdAHc+9y5hFwBhBQkbfwKhHCsb7rVeV9JJPYjtwDdLHosw
QsU2xSwJ7R4Bj1KimQq5PnX0ZtGVa9ReEptoV2ystE5kmX5K1Wpqtc2fs0CYvuk9
x9ZwnbLJ1CS27Az8LLoT36UauNJF2QtvUn6RCq0RbSMGMJsojvvKF48Rd84IfaNg
PPYLOahvp62eT16YIdRR4ob11G/L5zCqmfD2HqzNWV5UTvSiLIOe75LdkC1Bt+RQ
/35Tr9B0KETsAXMxvxaEMvBrfGPrsdc0cmssLyyGjGJkCuGVAq5LGu9WtH3rJQoU
qPo2VK2TqEfrtX40+tZFkNd8jMyUH588rD5sI3WY4aX+oE++EzP+gRMl/pTu6Rd7
jdwaJbInln43Lpxih4fOXEY3HlI2pqVGjsMg9mK2BOs6y7Tkqe/2S9MvjBCVz939
EwdKNw7b7rZGAZA+H/DV4JpaEFgeCzRc2OXGWhXQgpJlAXMO8KQiiqLzwuFrI+oZ
dkws0PhufR2JA7kfZKA5q2pwI0ysqDgJ2xPISao5tT6HAuy7rz2VM2isxX9/rpct
C2nsOqq7m0oNwPMhGBsfsT9Bj6wkVMZ6mBEyQLKFQNZmNeDw6l80ZobjeQaOnOGI
WBNwL1PLtfHcPQ6kfSNwyKHtmEh7Ap0PSKZ5YsPEdz4OHZ/XjbD8YFyJ451NuLmp
abFfYiMCmYy6tRFIy5XwmvL/4sUMPVzynjh/YQzdKMPY12on4PiTDmsABUTTkl32
Z/qGDkRt3BNHU56PoMLo9brFhhU/4MybjZO55u66UM/dN5E1nV0UQFTe7r9XHqDJ
jStSwIag+8g9w0L6S/kWEZgGj/MhZGuNFc4vGZKF8njk1MuvjZxhtYszi3YfUjwv
ggXZEqh5cPnITlmbDK+quVGsqWOQkRs6zetvOJEUAwV5KqBpzQZCB7el3sCXBDrE
sxGe0/Q5iUpj4Wmaz3W64rI+SSmOa9t2Mvi8+RF25GBwKXgpufho56fgSYwshOXG
AjA0qHWVycXx9nv0e8/fYPMAnl65wgaQV2ZiqdCMTI01cmV/jgekuD/pcf4nFV0O
CbkR8v5hMz8XR5ZKDMolv+8ySFiCPq0HsvyXNBJq0pFmS97y95w7dw6s5GLVJCnm
15kldBpnN/++hd2HSUXwF2FwfNDms+lCRUrf7KJs/GsxqrFUFB0fOGVQylxMA+w3
QDeVYTQ0JqR5xtsJZ8nu3I7hAxdzfb1XgM5pWYluMSj7PFVNrU0nxMWXrjBQ2tvf
zg3kgQB52aXTEKO1BUZHrNmepzaYdioGPdqpxQDye0aB0pqesXwwflWZ7/MbHNEg
PI8j3IQr5iScQSDF6pX3gWzmLxjE2q6pV9/Up/cbHN+SA5iQkETKQgiq8e5Bq0UX
468pkLFTuU60WlMrCKOZ6nIobPNsD9dVFdEWt5zfKRuUF6Etqt/KhLWfHV2w6YXn
C/rttBaSbUeC+aXZ+FcULWcj4Yb3CKyVwAHZ+ytugj4tEvG2Jz6aAKAfBtthUe6v
pxYG4toD6I7K+yhfRAMPgR7hrogB8Y6ilAhxl1Zh47nWqnjB3uGCGv0leMf0Ff0v
1zIMd2snHegOJfZZA9F4PG6POpgVZAOJJLHB/qtkTralbu5uDe1vpKbGPZPD9siX
dRPq5nBjJvUafcL8ZhQPILJTC+J/SdTl1zXSppF6XdixwxTbfQLRGO/hlvVj0MQx
GMsZmN90Lt545ih/Uk5tlSI4MHJ5ozM5dXkGP/+jyZ9TYuCfB5LxP9k43xwAcCzo
TwviBj7WNTSRttGI+/2tQRO8yRKr6mCpBPrikd7hU+LZ2irxa1n3D1W4XgI24pGo
qaOY0F8A9pk3BJDzUMZYl4nETnMPYxkHB3YA+boUTWTurB+Np64yWsUz7F1W8UYW
yL0q4Q0lrPrUV/iJLtSXE0xn+NAASQxWuTcaP+ZIciQfn9WE/O+g0/H+itJ+3Fgf
+rBPm5qs6N4o/4/QdDJZX2xNBmQ4W+OfKzBimzwLAOqmF1QmS2e1tW1ZniGxSXPe
DY+rQ3RxR/fboXmSH4YR7lJtS3/BR/KWx+Mu5LezWEwOwQGaviXDxZSDkfbDMbxw
+V2ZanQQv5fXEMZjsLQB8FKBpwW5KqHAq6Vgj5jQIeeJTAhJ8kw8/prbBxsTLACD
btbH0K81j7JzO8ibF0LLkfld/qtwjkAFg60TBvGikBXA7jrLp7f1HW/d10INZ6GR
RTOZEe386g5WYQqhKY+HTNa8BRpMejPkacNHU51t4Od7ntz6R4b6qqFvO9w+isH1
33n6ejEdWkzrI5M72w35+NPQ1+AQzmmwFRa1w2qLJS1ZfixTueSHQ8dvEip8+5K6
TE6531iq41PxUO0KJi43ixY4zsQf6ndnito0T9BgRn2cWr0re1DPCJ6NmcOGhjXZ
BH3SU5OyLhFK2pcjvsiaIQ281NI0FfSbZM8TUdGWc+wMO5HZrfB0LIdPZYagxwpN
N0qT5RukHUBQ2kl9HI0xRQjyk8IoXN2MihE+5TKFQ6wrBPxetcDlFo3+2/Phutcd
8WrhYO2jm7nnTj0K94HMPqbNHL62cnEpKeYb9UPyaouIWYbAJIfvZibvywjBnTwE
eK+PC7uXz+Ied1f2X3j08xA4I9cuvdFlHKlMJn8adc35ZHRf0IEgOml6F29T/+P9
tXb1KTHj86WYRwujzhu5tnFKSlra6EVQpDPnNo6iZAHRuLeSIdjErXNK6wpYoZmD
ak5Ztnm/d6i9E2NZENgncv5W1mcCqE4HWBSnGTuxIntQsaPTE1kYWBetYZ89o8H+
duSAVTOb3bvmkpZbT8huQEwc6bNmJsS06HPwTayzo6oLOX8Wg05Df9H6mo3a+Fgp
fc7WCg2xT+bmF0BRl2dalxjsj+8Q7GHXt8teRSyO69K2Z87X/PeyC3iLdGIavR5t
p4mpxUI51D7b7df1KNPFOJDSVP3/4MJbRs5QWY2zUUpWLCMk8GrBMhl4GE+/zLPZ
uujScJzHdFjTuj7tR6FTNS1+6V0xnoZBuaWqLkDL52/CHQS3tzhpjJfpinzWMRnG
FO+JWZ0RXaAz7XBU4nBnLcEiSuTvjmMITZ/mEKTvrDieB+chu5prYQwfEJ+hsRLB
Qm55bJAoYE30YaxHACBgzT3mbKMn6W+z9HZgsR/zrhqjuJck8CnjPPTIbRF5g0Zk
6mKf1xK95GW+t1y43XBFGIFI/5cLycv7vpFzT5YPK7fgoTfToO25j415qMTLVIm+
jCHCKW7jOonwiXUgi5MDwAyaQcJ1XrhrSGvolZAlGhcFH+sJ0wc+6mWMRjhuE69P
lWAhboS1r+f6G1Buzv7YneVrqDC6eCSy8ZJpG9AVaiGtjTSDSr/4X4Kaancoiq6u
bczVouOcH8YTXV0wi4h/uj9kPRCj0gu4nSI7yF8ooguVY3asbI/XtEdOPP2+Daga
jD+cmdBa8NBUxzWm9ZoTE0Mno2/uBU/P6P3zMsyspc7OLKuufab3u7qmiG7BRLeK
qLlOS+ao4qqmWKFFOCzTwmiOSzhokKsaMg5LDm4Z4e/k/fj+kcgzoztBsWrJmLyy
QANX38wpogLPt62GJW9Nc4qt5YyqilJYAvXd8hqHFRqM9LLBLVbkjMP4dce0az1u
5Jj6N04iWOCNphdnTCULAiwpXUvI9lw/6z6C2+1+tyeyflzK6XX6wwWycwKox0Q9
wpmGKmQCXkoAeuPnzPibYnZ8TlbL/Y32bPsoEWlDcSHMzrtnVFexMKEGTtt/lu9t
ifxXh4PpBYP+w+jYkwiG7rKAAczWyVXceyQyZEV3dGPfwptAQ26JnvPmv9/0k8M2
R0lfZHg+QS9tIyzCgeNi6ZoWoAAjZFXDuJBHkefGTY7W8vdj2BGBO2CuWA2g4FCH
yUZZ+k7gUNXlA2aUpfy7aTZB39pKHo9Eu1r/ZFXmiY607ExY9tII3PYsQJyKRUex
wJN2Rnnr3jCn//tvZKJPmJjPxJ/KxkZMW1dysMBTWnnbpcACK9WkDaNo9EkFMqL9
FyRwUTMaCQ/OcG7/ArJBPRrwPduhMJ6/Io4roni4o/mGTK+0/32nJ4erjjvDMJKW
QVLF6vr81yV6OIwX9LSzPTaS8cQx1dbloF3VRyHMSZ77RGAENlZ7SUOevcR5lLOJ
pVjiYxUvB+h3obwXWGjseSEBWPWeisKXCo8b/rO6p45AR/TRRv9rpokbsVRRDtPa
5NhlYiFJ3yM72hv1+NDZ/7KM5fAyAx5cabyoI5KzScxM/LtNWKIynH00zq3Epe5Q
SXbu48AGl6E9sQThRoCAHfXKpEPuF8GYiZmG+JfhvdX2HfjjKDKLnzWHmq+Eb5BP
cx83inF5zPKwrbO8NCPf6JTVorzK5L3uh2+h54c6fK/YjbnIXyhxQYvAlzY82C58
EgL5MyxWYs1uoYZ+ATStD13GOGLcMPSM5TZjQMcaWv86SV0gvMA7kPkgC7QfHjt3
cK/+v/f/F6XKV+am7rM6bnzifLMQZ+1zr3AtdFjjz/Vo/L27moFn6nZVVNrTBII1
+4D42QQTYCXbgoQ1HtwvzO5JKoZ/TxKb4Y7u+uxVzHFeaUYZuEnMzQUjZeNyX7V9
mEX6srks+7u9XGotms+jLDI8osUAyUl0CEg/E9TnY80XrqKFBEbbPYgkfGaGzRmN
+V+7qO9FJdkjNyM91mA/2HLoxgMz4X79utjwWSd7UYzdPtPY7B/nGusCUJUKHRwe
1Qa186fxBkzcBHCvfIsHaS4w3lC6+4NCkgRQu1AsOjRuZ+GN4hg4D27Nb09v9+rg
a9yTPXRLJVPJLAkgmMv/0PEGP6sOGI8DNAxN0a54LGSzTnguCBDSB4iZecyktFYT
31pSVKAPXPwcrvyW/jn6mXPY5kJAk4rCX+SC4auKsXmwo2AsxfUKfN+fTZ6vffis
2GqsktxEB0jKsllrf2zIVKr1nbWp2RhjX/SdFbxhoz9mkgSiRvDDgtz6lBan74ez
8egNBZxX5oBvnT5Sr9sQZt68SAFVxau+CuLE7ojgs26ff6ot9UDRt2dR0bq9Bzdu
xgOPLMwKe4Bh0FJtdI3/lrAHJ/N20HN3cswPOx/PZj61iw9LHPItTJLl8WLB8GaH
lUT6aUCQrtLmN8XK6BkuUKArF1FYkKPufBSGOiYFWh9MUmB4SgmJPEhd0DuiNaK4
WsiWe2qJA+oWfjKAPW93l5sALPpApHLEPT5qQ4O8gJ5s8mVM/U8jFgGXDH2lkmhM
jyVWVAIwr0O8e8g6p5iYhJA2MAJR2A1rnyz+LL4u4RDJGxRjHtlzUx4YYSDeoeRA
k2FtL2+7diqttUBEBtXXxT4o0kqn1QrXcOOY3kqaJU8VKMztE/wN01JOy/6pNG0c
THQrNPdVRXrPcQrOtc26eqOlhVlx9zQpHZD/PL+SusfhzQJj4YgpBrEB+HJh5IQV
8S87uSMgMaKIpFhDAWGn+agSl9s0tw0Z10zg23AZIlhMPmZCKbtZdzHUl05AdYhi
8/2sL92QuCdxHRRch/Q2K/Zxz2ClTpMeeilGeb7ImpKJ7/tseLHFrYwL0N3Spftn
OYziTjA1KIMQIcbVp3WvZXa9w36yQ0Y+EOl7U6MSNoB7dSGl7Ga3P3TjwP0i0irK
V6I7Htm5EDEJ1XgVxK6tUt47UhWrdTAKczfLfpLj8Vgwiyhxmbro1CHp758aKDAJ
afy2hMEt+BYP7TXmK8bmLKox8f5nU67oVD8+/CbsUIXRlQLvD2I2M89J03Ertyuo
BpZ6l+uOIjQbVAx88YQ2H1Ng4dvXZEatrOKd9lGd96Lvuz8l+52vRatQC5a8MMB8
GNPQlMjcvQQPJtSgmtmh2hSCcL/QN/lybiY0Dfg2QS+ZKYxvvKzs+RDLsci1WJUa
JHSlrLUjmOdbeRJDGGgzu/4DzLeDgWpO2sa7VoXEnvqHvBwQNccqC3BPnPG0kuG6
R4InMDtOgalq3sEathAJXlIrOKHWzTuSeDG36CktnhP2nBhAnNKAhQX9k3FGVudG
/erOFT7Vm4CSbZjCNK/zfdePwcnEVYurkqrVmJ1pVsXH+0oxbdFraMfCnWx8Ijo4
HcY/1HZ9M1S/lPXy0zmw+ugwD5ZuXDsZAvCBfuHsnPFu1T3lIP79+wy29BPTRRY/
gLvBskzhEIPy4eJ3vwshnBSOoWFSS1gbaFmO8RIhafAVdARhUKcLt95f9GuDJGLf
ze8YZE0HF6NNkMBSPvPFlt56kdQmsPR2WwNRBbYfOzrxSLicM8bygTIwqr1zl/dT
2Kbu+EYSLrEaNMdhcTkDmB984fKxfHsjBBJFK8Vn5nWhqRR7ubC0XS7pf/QbWa35
/vH1fwqU/gvAMvYAej7TWhT9nsvRbjCdpcVYDHcl3fECTYnQxjGNib3OxthM8FRQ
/nnAhpi/ObkhwIOh3XxyMlKC0eoj07Ou5XWj6LYLg2ag9/kDqysFKyPJCkC6KQa7
r5B9HxypIg5MtD+2GAsqMHlH0wyjeXGAYK57lWmdbHiByj0tiGo7+MNszQvh0rcZ
RZ+39A9k3qda/9BmnzuqBn/1ZeJo0TvFXZXG866uCXlxq3OvrgE58fcemY87d/q6
WoD0FEqntBJP72hYyvElwzLpwVnwImdFtEbz1l/QLiwxgoXOA8dDoNc/iVUFxnW8
aYA+5NrK1nHvY5gnmDq+eno//Oia6hqPF+HgRNsSpi3vm7uhyLsIsSEHkkW71IP1
BDsakKzYtFGrJpzPgFF1VxcfWee7UWzEHqMmiMIFa8jilKvKrIvKayISkky9nRmT
Lv07Wgreu96f+0Jsf2TRDWJpp6LXgz8OY7uBVCZk9x+iqXttrJCADs0Z7rNTn3cA
yUCCXD1UszBFEooRZrjB4h7FPojMDutAbDaLf+N1xQm9CzdJAob27tqjpNyR2Nme
WzZjuDY5Y+CuoAQJCY+A6N835VqvNqs2WLsM2OaTrK6MvRD/HvOLdq4TCMx4l51A
SdN92tFSQ/b/4n2PHf6m7npJip90FxD0QVK9dGHWUYStYUZz3d018Ileu1jMh9fk
e35Bp2nQ4sRaKASUCd6l/O+wc57YMcANT6JuPqZl1yS54lMKwHbWg0ZHkzjPfz6q
TnZGDo/7qEssSY6DccfLSjWbxGe3TypskiL7qK8tXqG+N0gMmm+3EoSWGXXJ6C70
1MaFTshU4fqMHB/hieDOtYBpTUAAAaetWyYCBiHfAg7AXOXZ56EItr0txfnlxhJW
3yhzEGZ1bpqMJ9/WgJC7fGWll1qo7+36/wJUfTl20E84GgeRbzB276dpm3/coyg9
nvwGxihnlpdV3L/f3ViAXC95XveOju/HqW7q1+JwckDneEsr5Y2SavXAJf8Ecgcy
mMxb7Sxk+sd2c9nPNpWBbhOBb4+J2i5ahoQKGHUsFFJYiGZpFpZIAa46J2vdR4Rk
Bwtr2Cyu3PyDT0of/BaitkJnbpoOy/VP3KTFv1JHX/mModWF5/V9C42kCpi6qR0G
8RgsoI4TyQhc4M8L6aO/KuwY8yU9Z2h4ZdrP/8DBQ8pQ5n+mn6boUudMFPBNOLlX
KmCWYbQ9EmnlWo6xcMNfdK/YxbKdCXplBH4wXFRmd2blGVFjpkVdQcZ1flOq9UjK
TVKzclsEVCo9v1PzRIR/4YPbxf1w4C41J0EDPd2O1to8EFwiOT/QfWETz6wIWF4j
Ii2AWlTWRcJFhqt9xsYKDvRr8FCuNZZ0eYjuQHRfcTNJQoOqjPjnjAPNoC2jQ6Hj
qQGqPy9rj3dW+pP3bf54uv07t2Ui/1Zlq5Qa8fcY1uOsl93wi7dliWdMyb0zmIzU
L7rdEybP8Al7LsNn/e/o3l98aEPDsdkU3LTM6BtPoVDTcfd4CmNiaTP9dRd9Zq63
l0Ez+Aq5kdapUEMG3E6h6KSarLyySEtuus9m+nOjDcnQDx/yPUBRnHKOlTSAG3Ox
sMTtxyidm3ruvn7PW9Yia3uUUjfy56Oe76fI1lTp9hZMnLFU4ic3/IDB+2P1yvUn
BSc1zB07YT0eAmyoLQN0nD83NcLXhO5w+67eUPG9NhzVwgvQDDslPfJLQYkLhjzS
CWH9HSePKcWJaBwZrW8MxDxi/QdXZ1UjcK9eF/O/Wp/Kb7tZbQ9ipnGjvDMgNzkf
9JIoJL3At5CQi0GnvRzHMnZZNCYCJ4vgOQgn02VyD6EjUNKDpOws/tnqmCIh1XTo
BQ/WgGcc0s5P4rmBnUPK8R8LH9kxCkbQqD7T93wyQeylboEbq9nw6A405rXUBQpl
u7qAPcwsKSEgYDrlIWydVhmMlzurmJ6RNId31Bqyo9xRyLD5YJuX0eex9b17MNDo
dVcGZueKzTHU8EwEALhO2KMj+Bb+Q4KwM8ZqL4YxgiBW5B1nwqhkxH+SCPT+ZNmp
yvPY0/UdNNeFd74exm2xrb2Ek/bzcANv3o5mYm9/O4nOYAtRwrkSuxzbbGxbc4R2
zdIISVJ2kACkwAZRZ0Y0Lm9FWj4M5VlHBMyTfi+66/hpvow2zEwNxO1+hMHJspj6
FLTmaffqNklMC3Y+t6gv1reRbQUn55b5PVQ0BLQZtT5zopr4Ip3yJHk81E3WU6tQ
Q/hk4Tt0/CXPrXsJu/3FaAucr7bjBDM/pJ1CBkIAK4MOU5Q/Xc3rM9ZgG/2U5kgh
IHMVZJ8lSEB1MMNQkBIDviuE1H5N1eWhtq7kBnic39+qgtIJHS8eaf9lmERmhhHg
xr4Tay5lr2hc8YPVDtYFfum5nTgjN8VcRFxO/snQMLWgsNTbISqcX/xCPxErYKXr
kJwFaTx/8Onch+Fp2v4b9hyBhWO5m6TL8oPoGPMrMyhFuwGxXwCmMdUk2luH7C7B
k3t7f7y537P5BQ10s/DvAJMAzCbywLMRSCWmxN8cASlp+V1uxod0N+l1eAVD9knQ
nEDWu2Q8xj0Q/oeDgcn3+ymfRZ24XdRpwCuOAmbhxYjp1TA7gRwKCtT3oV/kSQMI
qs4F+naNzCKVLhWzmwMq+tbXUydpCeyugZir8Oig7bybilFY5s9yPnPDXd9pElet
P5tfkfInpLnMxt1DqGekiEwGb/D3nqW3w759PMhXhf/VVXCv5bNED4kd2VI3xFzO
qQ8jpWZ+WIY09yv8yGoQurc4Cl1oFmhRcw1/J3PNXxrTerz/TIQdrV1dRkm4aDjA
c332QZAh4wMVxtPSNjt+ObZGTOuS0ixPBZ/XA5/8PpfrCiCjC3ebneVoemuV2MQI
TCwM2FKhKm26Tyx3APJjS+CeXw+678drQAQBHUNXueLg80IkxWa0FxHrNQ+Ew3Wq
nc67fCAY/QJeUkyAYyqPqJj7I28piaT+MHJuWmcuI2NvwaCagKk2yIiPeGI6YQtY
UesOrX+mJ0KGTXE4k1tfgVshU/gwSD82ehYAn3tuYEp4lbv6HJ9CL8//gbd3Qvsc
cHBDKhO3Dprh7BcnaKa7jLMOxBETBVF4uuEwFqiQzsbgBaYKgzG7Y0XT60u1e62o
m4rolI2y6A4+1zb6GdWmqR09mij8RD8maw4qCRy8XibuMmeX2Il6/2TASfJhGsi0
c/jG7A2evzCeZ19ornI2ifb+XawwUQQoWqLal/uecUKAAmAHlpOXX9u/Y3giCsKB
GQyknN1YZa5ao2z62LuUBU8lvLQECycow3I2v4yDcfUhybnFVncOjVHOgffF0egK
QHHJZOqibk8oDw6qRJbIsmQza8xjlulb0AVA5a3Qb42ekK0WoLOLl6n0o1Op26Qe
uZ+DSh/oU2Ptu7oTkpESEUoIWrp0mxD0b5sSMgczLOnj2olUb7uMOEwX1FNiVaGn
6+bRlCAST8LwZHdLBtJ/QahWabqg+o9dXb4o0vvCY68ypAwamey0o5Vt8gaa/s0n
oEVRc2x9G9iI3wxKMAMCLne1KfwaaNELrb3jxImzISflirYkPRdyYYaAX5O3YEic
ykqCK9Kx/q6zovA5dRG5ZmW6h1Ubf4aCFA8CJdp/g3ZDcE5tH8vpk903YSB+99zT
M3CVj+w9XXgjqKgZV2gA7h2FtCGIMCkRNjBV1RZfRcTyUoOb5w1Tse+J7ZLOLxGV
IhNxZRSqSVyIMcgWZTNMpG76sK74LLIBUs7pB1JR3G7j6l3peH9fjYEQgeMQuCcP
x1Df4nMWdUyEcZFtqbmVAsG+28kYij/JwPixHGQCJYLU+/uGh7gvFWkJGVXgTubp
G0CGUf1Tqv2tD1qcnPr8CVf2LyE5lxrKmUuF6FckXnEsnRKOt+w4TBf91kjSf2uF
oqKj2DCZ+4qD9cz2bANOty9r79wTuZT3VX/CUIrAVrJwuOHcUpeu2yC75hXuyvab
34WmDiM60Y+dm1tmJ3cuuTzby+YiUfEGf1s0SZJk0qypy2sjBhHMh7Ixo6YA+15P
qE4lDbIawnnUKbHw7ZPLgzKfdLYG/0uw7pRAk/mXjnU7GojhYvH8FkJgLulCOoml
tH5lVLY20cEi8mU8JuE1/NyM9W8/k34Tl9TUFZ0hqUw0Pzfu6MJ939aUqKVl7huj
R6H108O6e8jVllIyJA0f0Mlg8L0jaFvLQ0GlDeaYIKDBq6wri9UC9tDlPh2zNtBq
YugLUIUaiSztmnSfwE3tS8tlrK/YORG1aoKheqLdJTrP9QgJn84YxrLCEbcNc8M7
iGcJ1PCpDMJKtvOF94buQoqDP+SJP6tNg64F1OzF/2J9WFr8Vrp2proovTD74IQo
m1vTci5HKW1yAVNLAK7kj++O95Y6Qw8Ehn3NPgcljPgFquZcBJbIE7YWw84YvRNK
kXNYfch9Z9jnNuW2iJZ8Blbl1iViBejNoQKgF89V03TDIELXOL66ZVnIK2bNSyuX
QmCYLJNEvo/GZuCYKXz/V8h+PswcbaOKMET0sr+Z5o/IVVmruIwS7qdxpzKA9G/C
fmmJPREXI1YMnipvDfnCYqbKgMZhQD7lkX7VlacNkdw839orTuGV7gbCljBOBAud
Je/aSu29y4GeAm+dVKE/V613g32OoH+F/Lrh65kHSdYbTtv/6CMF7gNvT4MIVRJD
8rHxr1e+DrouobBDefrA0b8BQOWr/3ArPO3+QtjCW2iEf27t/I0JIm9P2dyb/p+4
6pmdt4jc86PTNXXq3HsDKSV0fnPNezIx4RIhmEIVXW6+Fhwvln2/le6/+6eg0m/O
Ti3cGgKwbMNccfk/EDNR8vGk955M3B5NpguOv4ZeXmA8VbcXHSdJvUdqL4CFtmtS
oDi/SQviltOnVaEbBkiHpw/R9yTlXgYD+O8xT/DwdF5hKIo7PHB6mKjbx+K6XsGu
aqwX8y8H/6k06JAeeXdTLLiO/CLx+tzrt4Ryiyn2EXFoaW11sBHrF3lLaRpiNR8G
XFkroDlceS0iCb+z67Ge/3LqVrbtpoB7Z203gtCsWJoEBHfULDdHzvU+0CBuSzEw
m0xkP5J3140rPcSeCX1GK1pEEQYUr17yEDomVnJoQ/33MRgUW1yY3QYa3xGvQ4Nb
C2UvqncfyrzTeCfbPVhbCH5GOJk62oYbv0vh2SdurmVoJ8lgBSi1pzvOH2syHkWP
UXk+hxswFI7jv29e9pGUAh5EBTpQLgJkuwLCy8dk1n0R1XtUVBirxjh8wVZDJhPG
/UpP8LZF5Gu1Cp9jKhRCTQ==
`pragma protect end_protected
