// megafunction wizard: %Jesd204b v14.0%
// GENERATION: XML
// altera_jesd204.v

// Generated using ACDS version 14.0 200 at 2014.07.17.13:20:13

`timescale 1 ps / 1 ps
module altera_jesd204 (
		input  wire         tx_pll_ref_clk,             //            tx_pll_ref_clk.clk
		input  wire         txlink_clk,                 //                txlink_clk.clk
		input  wire         txlink_rst_n_reset_n,       //              txlink_rst_n.reset_n
		input  wire         jesd204_tx_avs_clk,         //        jesd204_tx_avs_clk.clk
		input  wire         jesd204_tx_avs_rst_n,       //      jesd204_tx_avs_rst_n.reset_n
		input  wire         jesd204_tx_avs_chipselect,  //            jesd204_tx_avs.chipselect
		input  wire [7:0]   jesd204_tx_avs_address,     //                          .address
		input  wire         jesd204_tx_avs_read,        //                          .read
		output wire [31:0]  jesd204_tx_avs_readdata,    //                          .readdata
		output wire         jesd204_tx_avs_waitrequest, //                          .waitrequest
		input  wire         jesd204_tx_avs_write,       //                          .write
		input  wire [31:0]  jesd204_tx_avs_writedata,   //                          .writedata
		input  wire [63:0]  jesd204_tx_link_data,       //           jesd204_tx_link.data
		input  wire         jesd204_tx_link_valid,      //                          .valid
		output wire         jesd204_tx_link_ready,      //                          .ready
		output wire         jesd204_tx_int,             //            jesd204_tx_int.export
		input  wire         tx_sysref,                  //                 tx_sysref.export
		input  wire         sync_n,                     //                    sync_n.export
		output wire         tx_dev_sync_n,              //             tx_dev_sync_n.export
		input  wire         mdev_sync_n,                //               mdev_sync_n.export
		output wire         jesd204_tx_frame_ready,     //    jesd204_tx_frame_ready.export
		output wire [4:0]   tx_csr_l,                   //                  tx_csr_l.export
		output wire [7:0]   tx_csr_f,                   //                  tx_csr_f.export
		output wire [4:0]   tx_csr_k,                   //                  tx_csr_k.export
		output wire [7:0]   tx_csr_m,                   //                  tx_csr_m.export
		output wire [1:0]   tx_csr_cs,                  //                 tx_csr_cs.export
		output wire [4:0]   tx_csr_n,                   //                  tx_csr_n.export
		output wire [4:0]   tx_csr_np,                  //                 tx_csr_np.export
		output wire [4:0]   tx_csr_s,                   //                  tx_csr_s.export
		output wire         tx_csr_hd,                  //                 tx_csr_hd.export
		output wire [4:0]   tx_csr_cf,                  //                 tx_csr_cf.export
		output wire [1:0]   tx_csr_lane_powerdown,      //     tx_csr_lane_powerdown.export
		output wire [3:0]   csr_tx_testmode,            //           csr_tx_testmode.export
		output wire [31:0]  csr_tx_testpattern_a,       //      csr_tx_testpattern_a.export
		output wire [31:0]  csr_tx_testpattern_b,       //      csr_tx_testpattern_b.export
		output wire [31:0]  csr_tx_testpattern_c,       //      csr_tx_testpattern_c.export
		output wire [31:0]  csr_tx_testpattern_d,       //      csr_tx_testpattern_d.export
		input  wire         jesd204_tx_frame_error,     //    jesd204_tx_frame_error.export
		output wire [63:0]  jesd204_tx_dlb_data,        //       jesd204_tx_dlb_data.export
		output wire [7:0]   jesd204_tx_dlb_kchar_data,  // jesd204_tx_dlb_kchar_data.export
		output wire [1:0]   txphy_clk,                  //                 txphy_clk.tx_std_clkout
		output wire [1:0]   tx_serial_data,             //            tx_serial_data.tx_serial_data
		input  wire [0:0]   pll_powerdown,              //             pll_powerdown.pll_powerdown
		input  wire [1:0]   tx_analogreset,             //            tx_analogreset.tx_analogreset
		input  wire [1:0]   tx_digitalreset,            //           tx_digitalreset.tx_digitalreset
		output wire [1:0]   pll_locked,                 //                pll_locked.export
		output wire [1:0]   tx_cal_busy,                //               tx_cal_busy.export
		input  wire         rx_pll_ref_clk,             //            rx_pll_ref_clk.clk
		input  wire         rxlink_clk,                 //                rxlink_clk.clk
		input  wire         rxlink_rst_n_reset_n,       //              rxlink_rst_n.reset_n
		input  wire         jesd204_rx_avs_clk,         //        jesd204_rx_avs_clk.clk
		input  wire         jesd204_rx_avs_rst_n,       //      jesd204_rx_avs_rst_n.reset_n
		input  wire         jesd204_rx_avs_chipselect,  //            jesd204_rx_avs.chipselect
		input  wire [7:0]   jesd204_rx_avs_address,     //                          .address
		input  wire         jesd204_rx_avs_read,        //                          .read
		output wire [31:0]  jesd204_rx_avs_readdata,    //                          .readdata
		output wire         jesd204_rx_avs_waitrequest, //                          .waitrequest
		input  wire         jesd204_rx_avs_write,       //                          .write
		input  wire [31:0]  jesd204_rx_avs_writedata,   //                          .writedata
		output wire [63:0]  jesd204_rx_link_data,       //           jesd204_rx_link.data
		output wire         jesd204_rx_link_valid,      //                          .valid
		input  wire         jesd204_rx_link_ready,      //                          .ready
		input  wire [63:0]  jesd204_rx_dlb_data,        //       jesd204_rx_dlb_data.export
		input  wire [1:0]   jesd204_rx_dlb_data_valid,  // jesd204_rx_dlb_data_valid.export
		input  wire [7:0]   jesd204_rx_dlb_kchar_data,  // jesd204_rx_dlb_kchar_data.export
		input  wire [7:0]   jesd204_rx_dlb_errdetect,   //  jesd204_rx_dlb_errdetect.export
		input  wire [7:0]   jesd204_rx_dlb_disperr,     //    jesd204_rx_dlb_disperr.export
		input  wire         alldev_lane_aligned,        //       alldev_lane_aligned.export
		input  wire         rx_sysref,                  //                 rx_sysref.export
		input  wire         jesd204_rx_frame_error,     //    jesd204_rx_frame_error.export
		output wire         jesd204_rx_int,             //            jesd204_rx_int.export
		output wire [3:0]   csr_rx_testmode,            //           csr_rx_testmode.export
		output wire         dev_lane_aligned,           //          dev_lane_aligned.export
		output wire         rx_dev_sync_n,              //             rx_dev_sync_n.export
		output wire [3:0]   rx_sof,                     //                    rx_sof.export
		output wire [3:0]   rx_somf,                    //                   rx_somf.export
		output wire [7:0]   rx_csr_f,                   //                  rx_csr_f.export
		output wire [4:0]   rx_csr_k,                   //                  rx_csr_k.export
		output wire [4:0]   rx_csr_l,                   //                  rx_csr_l.export
		output wire [7:0]   rx_csr_m,                   //                  rx_csr_m.export
		output wire [4:0]   rx_csr_n,                   //                  rx_csr_n.export
		output wire [4:0]   rx_csr_s,                   //                  rx_csr_s.export
		output wire [4:0]   rx_csr_cf,                  //                 rx_csr_cf.export
		output wire [1:0]   rx_csr_cs,                  //                 rx_csr_cs.export
		output wire         rx_csr_hd,                  //                 rx_csr_hd.export
		output wire [4:0]   rx_csr_np,                  //                 rx_csr_np.export
		output wire [1:0]   rx_csr_lane_powerdown,      //     rx_csr_lane_powerdown.export
		output wire [1:0]   rxphy_clk,                  //                 rxphy_clk.rx_std_clkout
		input  wire [1:0]   rx_serial_data,             //            rx_serial_data.rx_serial_data
		input  wire [1:0]   rx_analogreset,             //            rx_analogreset.rx_analogreset
		input  wire [1:0]   rx_digitalreset,            //           rx_digitalreset.rx_digitalreset
		input  wire [209:0] reconfig_to_xcvr,           //          reconfig_to_xcvr.reconfig_to_xcvr
		output wire [137:0] reconfig_from_xcvr,         //        reconfig_from_xcvr.reconfig_from_xcvr
		output wire [1:0]   rx_islockedtodata,          //         rx_islockedtodata.export
		output wire [1:0]   rx_cal_busy,                //               rx_cal_busy.export
		input  wire [1:0]   rx_seriallpbken             //           rx_seriallpbken.rx_seriallpbken
	);

	altera_jesd204_0002 #(
		.DEVICE_FAMILY            ("Arria V"),
		.SUBCLASSV                (1),
		.PCS_CONFIG               ("JESD_PCS_CFG1"),
		.L                        (2),
		.M                        (2),
		.F                        (2),
		.N                        (14),
		.N_PRIME                  (16),
		.S                        (1),
		.K                        (32),
		.SCR                      (1),
		.CS                       (0),
		.CF                       (0),
		.HD                       (0),
		.ECC_EN                   (1),
		.DLB_TEST                 (0),
		.PHADJ                    (0),
		.ADJCNT                   (0),
		.ADJDIR                   (0),
		.OPTIMIZE                 (0),
		.DID                      (0),
		.BID                      (0),
		.LID0                     (0),
		.FCHK0                    (65),
		.LID1                     (1),
		.FCHK1                    (66),
		.LID2                     (2),
		.FCHK2                    (0),
		.LID3                     (3),
		.FCHK3                    (0),
		.LID4                     (4),
		.FCHK4                    (0),
		.LID5                     (5),
		.FCHK5                    (0),
		.LID6                     (6),
		.FCHK6                    (0),
		.LID7                     (7),
		.FCHK7                    (0),
		.JESDV                    (1),
		.PMA_WIDTH                (32),
		.SER_SIZE                 (4),
		.FK                       (64),
		.RES1                     (0),
		.RES2                     (0),
		.BIT_REVERSAL             (0),
		.BYTE_REVERSAL            (0),
		.ALIGNMENT_PATTERN        (658812),
		.PULSE_WIDTH              (2),
		.LS_FIFO_DEPTH            (32),
		.LS_FIFO_WIDTHU           (5),
		.UNUSED_TX_PARALLEL_WIDTH (8),
		.UNUSED_RX_PARALLEL_WIDTH (8),
		.XCVR_PLL_LOCKED_WIDTH    (1)
	) altera_jesd204_inst (
		.tx_pll_ref_clk             (tx_pll_ref_clk),             //            tx_pll_ref_clk.clk
		.txlink_clk                 (txlink_clk),                 //                txlink_clk.clk
		.txlink_rst_n_reset_n       (txlink_rst_n_reset_n),       //              txlink_rst_n.reset_n
		.jesd204_tx_avs_clk         (jesd204_tx_avs_clk),         //        jesd204_tx_avs_clk.clk
		.jesd204_tx_avs_rst_n       (jesd204_tx_avs_rst_n),       //      jesd204_tx_avs_rst_n.reset_n
		.jesd204_tx_avs_chipselect  (jesd204_tx_avs_chipselect),  //            jesd204_tx_avs.chipselect
		.jesd204_tx_avs_address     (jesd204_tx_avs_address),     //                          .address
		.jesd204_tx_avs_read        (jesd204_tx_avs_read),        //                          .read
		.jesd204_tx_avs_readdata    (jesd204_tx_avs_readdata),    //                          .readdata
		.jesd204_tx_avs_waitrequest (jesd204_tx_avs_waitrequest), //                          .waitrequest
		.jesd204_tx_avs_write       (jesd204_tx_avs_write),       //                          .write
		.jesd204_tx_avs_writedata   (jesd204_tx_avs_writedata),   //                          .writedata
		.jesd204_tx_link_data       (jesd204_tx_link_data),       //           jesd204_tx_link.data
		.jesd204_tx_link_valid      (jesd204_tx_link_valid),      //                          .valid
		.jesd204_tx_link_ready      (jesd204_tx_link_ready),      //                          .ready
		.jesd204_tx_int             (jesd204_tx_int),             //            jesd204_tx_int.export
		.tx_sysref                  (tx_sysref),                  //                 tx_sysref.export
		.sync_n                     (sync_n),                     //                    sync_n.export
		.tx_dev_sync_n              (tx_dev_sync_n),              //             tx_dev_sync_n.export
		.mdev_sync_n                (mdev_sync_n),                //               mdev_sync_n.export
		.jesd204_tx_frame_ready     (jesd204_tx_frame_ready),     //    jesd204_tx_frame_ready.export
		.tx_csr_l                   (tx_csr_l),                   //                  tx_csr_l.export
		.tx_csr_f                   (tx_csr_f),                   //                  tx_csr_f.export
		.tx_csr_k                   (tx_csr_k),                   //                  tx_csr_k.export
		.tx_csr_m                   (tx_csr_m),                   //                  tx_csr_m.export
		.tx_csr_cs                  (tx_csr_cs),                  //                 tx_csr_cs.export
		.tx_csr_n                   (tx_csr_n),                   //                  tx_csr_n.export
		.tx_csr_np                  (tx_csr_np),                  //                 tx_csr_np.export
		.tx_csr_s                   (tx_csr_s),                   //                  tx_csr_s.export
		.tx_csr_hd                  (tx_csr_hd),                  //                 tx_csr_hd.export
		.tx_csr_cf                  (tx_csr_cf),                  //                 tx_csr_cf.export
		.tx_csr_lane_powerdown      (tx_csr_lane_powerdown),      //     tx_csr_lane_powerdown.export
		.csr_tx_testmode            (csr_tx_testmode),            //           csr_tx_testmode.export
		.csr_tx_testpattern_a       (csr_tx_testpattern_a),       //      csr_tx_testpattern_a.export
		.csr_tx_testpattern_b       (csr_tx_testpattern_b),       //      csr_tx_testpattern_b.export
		.csr_tx_testpattern_c       (csr_tx_testpattern_c),       //      csr_tx_testpattern_c.export
		.csr_tx_testpattern_d       (csr_tx_testpattern_d),       //      csr_tx_testpattern_d.export
		.jesd204_tx_frame_error     (jesd204_tx_frame_error),     //    jesd204_tx_frame_error.export
		.jesd204_tx_dlb_data        (jesd204_tx_dlb_data),        //       jesd204_tx_dlb_data.export
		.jesd204_tx_dlb_kchar_data  (jesd204_tx_dlb_kchar_data),  // jesd204_tx_dlb_kchar_data.export
		.txphy_clk                  (txphy_clk),                  //                 txphy_clk.tx_std_clkout
		.tx_serial_data             (tx_serial_data),             //            tx_serial_data.tx_serial_data
		.pll_powerdown              (pll_powerdown),              //             pll_powerdown.pll_powerdown
		.tx_analogreset             (tx_analogreset),             //            tx_analogreset.tx_analogreset
		.tx_digitalreset            (tx_digitalreset),            //           tx_digitalreset.tx_digitalreset
		.pll_locked                 (pll_locked),                 //                pll_locked.export
		.tx_cal_busy                (tx_cal_busy),                //               tx_cal_busy.export
		.rx_pll_ref_clk             (rx_pll_ref_clk),             //            rx_pll_ref_clk.clk
		.rxlink_clk                 (rxlink_clk),                 //                rxlink_clk.clk
		.rxlink_rst_n_reset_n       (rxlink_rst_n_reset_n),       //              rxlink_rst_n.reset_n
		.jesd204_rx_avs_clk         (jesd204_rx_avs_clk),         //        jesd204_rx_avs_clk.clk
		.jesd204_rx_avs_rst_n       (jesd204_rx_avs_rst_n),       //      jesd204_rx_avs_rst_n.reset_n
		.jesd204_rx_avs_chipselect  (jesd204_rx_avs_chipselect),  //            jesd204_rx_avs.chipselect
		.jesd204_rx_avs_address     (jesd204_rx_avs_address),     //                          .address
		.jesd204_rx_avs_read        (jesd204_rx_avs_read),        //                          .read
		.jesd204_rx_avs_readdata    (jesd204_rx_avs_readdata),    //                          .readdata
		.jesd204_rx_avs_waitrequest (jesd204_rx_avs_waitrequest), //                          .waitrequest
		.jesd204_rx_avs_write       (jesd204_rx_avs_write),       //                          .write
		.jesd204_rx_avs_writedata   (jesd204_rx_avs_writedata),   //                          .writedata
		.jesd204_rx_link_data       (jesd204_rx_link_data),       //           jesd204_rx_link.data
		.jesd204_rx_link_valid      (jesd204_rx_link_valid),      //                          .valid
		.jesd204_rx_link_ready      (jesd204_rx_link_ready),      //                          .ready
		.jesd204_rx_dlb_data        (jesd204_rx_dlb_data),        //       jesd204_rx_dlb_data.export
		.jesd204_rx_dlb_data_valid  (jesd204_rx_dlb_data_valid),  // jesd204_rx_dlb_data_valid.export
		.jesd204_rx_dlb_kchar_data  (jesd204_rx_dlb_kchar_data),  // jesd204_rx_dlb_kchar_data.export
		.jesd204_rx_dlb_errdetect   (jesd204_rx_dlb_errdetect),   //  jesd204_rx_dlb_errdetect.export
		.jesd204_rx_dlb_disperr     (jesd204_rx_dlb_disperr),     //    jesd204_rx_dlb_disperr.export
		.alldev_lane_aligned        (alldev_lane_aligned),        //       alldev_lane_aligned.export
		.rx_sysref                  (rx_sysref),                  //                 rx_sysref.export
		.jesd204_rx_frame_error     (jesd204_rx_frame_error),     //    jesd204_rx_frame_error.export
		.jesd204_rx_int             (jesd204_rx_int),             //            jesd204_rx_int.export
		.csr_rx_testmode            (csr_rx_testmode),            //           csr_rx_testmode.export
		.dev_lane_aligned           (dev_lane_aligned),           //          dev_lane_aligned.export
		.rx_dev_sync_n              (rx_dev_sync_n),              //             rx_dev_sync_n.export
		.rx_sof                     (rx_sof),                     //                    rx_sof.export
		.rx_somf                    (rx_somf),                    //                   rx_somf.export
		.rx_csr_f                   (rx_csr_f),                   //                  rx_csr_f.export
		.rx_csr_k                   (rx_csr_k),                   //                  rx_csr_k.export
		.rx_csr_l                   (rx_csr_l),                   //                  rx_csr_l.export
		.rx_csr_m                   (rx_csr_m),                   //                  rx_csr_m.export
		.rx_csr_n                   (rx_csr_n),                   //                  rx_csr_n.export
		.rx_csr_s                   (rx_csr_s),                   //                  rx_csr_s.export
		.rx_csr_cf                  (rx_csr_cf),                  //                 rx_csr_cf.export
		.rx_csr_cs                  (rx_csr_cs),                  //                 rx_csr_cs.export
		.rx_csr_hd                  (rx_csr_hd),                  //                 rx_csr_hd.export
		.rx_csr_np                  (rx_csr_np),                  //                 rx_csr_np.export
		.rx_csr_lane_powerdown      (rx_csr_lane_powerdown),      //     rx_csr_lane_powerdown.export
		.rxphy_clk                  (rxphy_clk),                  //                 rxphy_clk.rx_std_clkout
		.rx_serial_data             (rx_serial_data),             //            rx_serial_data.rx_serial_data
		.rx_analogreset             (rx_analogreset),             //            rx_analogreset.rx_analogreset
		.rx_digitalreset            (rx_digitalreset),            //           rx_digitalreset.rx_digitalreset
		.reconfig_to_xcvr           (reconfig_to_xcvr),           //          reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr         (reconfig_from_xcvr),         //        reconfig_from_xcvr.reconfig_from_xcvr
		.rx_islockedtodata          (rx_islockedtodata),          //         rx_islockedtodata.export
		.rx_cal_busy                (rx_cal_busy),                //               rx_cal_busy.export
		.rx_seriallpbken            (rx_seriallpbken)             //           rx_seriallpbken.rx_seriallpbken
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2014 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_jesd204" version="14.0" >
// Retrieval info: 	<generic name="wrapper_opt" value="base_phy" />
// Retrieval info: 	<generic name="sdc_constraint" value="1.0" />
// Retrieval info: 	<generic name="DEVICE_FAMILY" value="Arria V" />
// Retrieval info: 	<generic name="DATA_PATH" value="RX_TX" />
// Retrieval info: 	<generic name="SUBCLASSV" value="1" />
// Retrieval info: 	<generic name="lane_rate" value="4915.0" />
// Retrieval info: 	<generic name="PCS_CONFIG" value="JESD_PCS_CFG1" />
// Retrieval info: 	<generic name="pll_type" value="CMU" />
// Retrieval info: 	<generic name="bonded_mode" value="bonded" />
// Retrieval info: 	<generic name="REFCLK_FREQ" value="122.875" />
// Retrieval info: 	<generic name="pll_reconfig_enable" value="false" />
// Retrieval info: 	<generic name="bitrev_en" value="false" />
// Retrieval info: 	<generic name="L" value="2" />
// Retrieval info: 	<generic name="M" value="2" />
// Retrieval info: 	<generic name="N" value="14" />
// Retrieval info: 	<generic name="N_PRIME" value="16" />
// Retrieval info: 	<generic name="S" value="1" />
// Retrieval info: 	<generic name="K" value="32" />
// Retrieval info: 	<generic name="SCR" value="1" />
// Retrieval info: 	<generic name="CS" value="0" />
// Retrieval info: 	<generic name="CF" value="0" />
// Retrieval info: 	<generic name="HD" value="0" />
// Retrieval info: 	<generic name="ECC_EN" value="1" />
// Retrieval info: 	<generic name="DLB_TEST" value="0" />
// Retrieval info: 	<generic name="PHADJ" value="0" />
// Retrieval info: 	<generic name="ADJCNT" value="0" />
// Retrieval info: 	<generic name="ADJDIR" value="0" />
// Retrieval info: 	<generic name="OPTIMIZE" value="0" />
// Retrieval info: 	<generic name="DID" value="0" />
// Retrieval info: 	<generic name="BID" value="0" />
// Retrieval info: 	<generic name="LID0" value="0" />
// Retrieval info: 	<generic name="LID1" value="1" />
// Retrieval info: 	<generic name="LID2" value="2" />
// Retrieval info: 	<generic name="LID3" value="3" />
// Retrieval info: 	<generic name="LID4" value="4" />
// Retrieval info: 	<generic name="LID5" value="5" />
// Retrieval info: 	<generic name="LID6" value="6" />
// Retrieval info: 	<generic name="LID7" value="7" />
// Retrieval info: 	<generic name="JESDV" value="1" />
// Retrieval info: 	<generic name="RES1" value="0" />
// Retrieval info: 	<generic name="RES2" value="0" />
// Retrieval info: 	<generic name="TEST_COMPONENTS_EN" value="false" />
// Retrieval info: 	<generic name="TERMINATE_RECONFIG_EN" value="false" />
// Retrieval info: 	<generic name="AUTO_DEVICE" value="Unknown" />
// Retrieval info: </instance>
// IPFS_FILES : altera_jesd204.vo
// RELATED_FILES: altera_jesd204.v, altera_jesd204_0002.v, altera_jesd204_rx_base.v, altera_jesd204_rx_csr.v, altera_jesd204_rx_ctl.v, altera_jesd204_rx_descrambler.v, altera_jesd204_rx_dll.v, altera_jesd204_rx_dll_char_val.v, altera_jesd204_rx_dll_cs.v, altera_jesd204_rx_dll_fs_char_replace.v, altera_jesd204_rx_dll_frame_align.v, altera_jesd204_rx_dll_lane_align.v, altera_jesd204_rx_dll_data_store.v, altera_jesd204_rx_dll_ecc_enc.v, altera_jesd204_rx_dll_ecc_dec.v, altera_jesd204_rx_dll_ecc_fifo.v, altera_jesd204_rx_dll_wo_ecc_fifo.v, altera_jesd204_rx_regmap.v, altera_jesd204_tx_base.v, altera_jesd204_tx_csr.v, altera_jesd204_tx_ctl.v, altera_jesd204_tx_dll.v, altera_jesd204_tx_regmap.v, altera_jesd204_tx_regmap_opt.v, altera_jesd204_tx_scrambler.v, altera_jesd204_inst_phy.v, altera_jesd204_tx_mlpcs.v, altera_jesd204_8b10b_enc.v, altera_jesd204_tx_pcs.v, altera_jesd204_wys_lut.v, altera_jesd204_xn_8b10b_enc.v, altera_jesd204_rx_mlpcs.v, altera_jesd204_8b10b_dec.v, altera_jesd204_rx_pcs.v, altera_jesd204_wa.v, altera_jesd204_xn_8b10b_dec.v, altera_jesd204_phy_adapter.v, altera_xcvr_functions.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, av_xcvr_h.sv, av_xcvr_avmm_csr.sv, av_tx_pma_ch.sv, av_tx_pma.sv, av_rx_pma.sv, av_pma.sv, av_pcs_ch.sv, av_pcs.sv, av_xcvr_avmm.sv, av_xcvr_native.sv, av_xcvr_plls.sv, av_xcvr_data_adapter.sv, av_reconfig_bundle_to_basic.sv, av_reconfig_bundle_to_xcvr.sv, av_hssi_8g_rx_pcs_rbc.sv, av_hssi_8g_tx_pcs_rbc.sv, av_hssi_common_pcs_pma_interface_rbc.sv, av_hssi_common_pld_pcs_interface_rbc.sv, av_hssi_pipe_gen1_2_rbc.sv, av_hssi_rx_pcs_pma_interface_rbc.sv, av_hssi_rx_pld_pcs_interface_rbc.sv, av_hssi_tx_pcs_pma_interface_rbc.sv, av_hssi_tx_pld_pcs_interface_rbc.sv, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_xcvr_native_av_functions_h.sv, altera_xcvr_native_av.sv, altera_xcvr_data_adapter_av.sv
