// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
O4mFlsDIFRbVpSTwS7UR/IGhbqfmdR3aXQSGkgG1RfY2BhWsCJmgTik+BNc4WEBn
2ZCStV5T7AAGtdVGhh+FJ+Vpv7cIHYQCAgHRQIpyA48RRAzqWolgHUuDYEXEQKlH
DrcxaAI/Fu6VtmvUIV4iIV9lg/P29BPYBepT2hr09wo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1856)
9jUYkdgCFRIRwm3kJrEBRhjY7mkxbg2L8ANsFq1lwJ/MBO4qG47ks0ovwKukp198
QiLuy5e+fF6WbEBueFtRwvvgafaKrsJGOP+ePWkfa764PcHFsoFGsQCj93CXV3EH
Jxsd8lhsux7AApj7VE170O0FBlTXKAtxNgmzs0ApnbwoUl0lpNMoISnXjgzWD8Om
ZOcAsZkAX0nxeX/eS0csBkxxAVWscBclBUPda4GLyha+Xeag6aZoETVKmSF3vGjW
PMSIZ9oxehuWHK5OWxJN4hwFMPXmNApaIOlF32v80cJgnpIkOdbR2MWifsz/E4p6
4YXD/xUDoe9JSPziVLqbWqnO30oXL6jtGqqcULk6Gtv37BEbXvcZoiAjfP1P7Jvf
aTqTelgje4YslnnNnIJHLSqAPDqx4xQcotvnCW+o+IXMwa8N9Kz6F/TF3KPY9BNd
Xu2ireoo89TvWmuRUUWeAxV2BoeswCfMFq2kGcBcxGpNpsTfLDkccGlgSr5dEogX
ZCttpYPTWKYZXdWk8o2viFi+IppzJJ0+xZjYnSxEvdCsG79AIQxBUX9EqFkYNPiy
WmxDT/7PQ9xsgDcgWcex8Sy0xgkSHY4JXxUhDHAiyXAoySjDJCUE7KLJT7kEDxuW
DYrwk03RDtkIdfMSE5ResF1RH/jp+GR/BkcEqgcMEwtu3xc/DhQrq8gv+ygeg/L7
7FR21iQeCCUtFbVzMJZiafGsepDHTr0fpaW9Z1WsAq+WYbnB31mfoGbV1Jb0XwKG
0AUtLBmXSalVrkk6HYxAZJlUZiYbVF6iucXzY3DHiLoJRqnXI6wEkxJepKjTnp7+
cA+FnJyYFkKyfqr5+s/IDewvx1DdqTn6EMBa+MGOjY3JlVTirm+aDPXWKtPzmeju
PZ3kiXchsfp4ZKEobcsxeL3UeV1hHHSt1Br3+4lwYNnp0Xlh5HBTp6KjkZeisyBs
Y+35o1BtFE4L+bxx2cmNP70deouDWl1sZF+nSk19Ag2mdfosMz+kPwn/pYwLf17T
WSYuovmCR+/W98eXWolaFOVFdIkU8YRPxkR4T1wcJVvzRSCnWywppl8YYqREr83u
0e/z6PhFPgbXuePtkTNHHxDehB3+CKB2WupeVTALz41G3AbMKsOJO4nfY+/i1a3q
8UuLmQjU/wP+H7vavp/FHIgKyWlSEfTUWW9BBHm3Hjzsx4KqXor5oAmpLibnCj1D
CSNuXuq+wLRszD0nQ0F41jrufXpbLfYopXrcS9abBD/PtGHf9o1I1cQwokasm9fv
XeQkjtXCvyBzGNAJcQnbpXYEFu0WmxNh4qKIF67q2SP1QUX9iSfFMMMQ0DN3AZTz
3Bx4dBHrQh4f2LJzDX/zK70KgV7vxrt1a0Y/tuIo7aYb5EncOvDHNHnoIYyHIaHS
gvujE6ybUE2LKqHusW6wb4efgJ+KRw2rSrY3qN5oddPahb/+zGU8gmyiAAp5Ftk3
qv3w+6XdKZWC7FUae48m6jgEOe6jZs6IdzA+30rGwEzNc4ho0gBuYEWC9/ykBi51
HBDJVzf6hTlJlBBPTyFenQ4yylVG7UA2K96HPSFnQadtpprO9/ZjGNLdOlN4Kpos
ttfOF6QOhbA26BUwjOwtRBlILoCBFzXcNQV98Fny4TRvUhz2ro6kXuePnI3x6L9f
H/ZRezgWCqZmTJlKtHPs+6TdhDXkLcdEDTcMo8KSihA9wlqM0RVZ8mY1xJgTYiPb
zO3pZ2hgeHoBoh1wdEWtui8EZ+U8R+YOfJlKkP1XEc3iAVjZ++6cfilpmvW48q3g
q1uYbDz6KwxRrIYcqUHICeVdujzgxxdxfzSjK/9UpdgW3y6SctUqqq/o60tTEvoH
iVLFKfxKPgUxn50d3GBSUGiWngORF/Es7V3+kP5shgBMoFxWzIQaS9qij96fyS05
3T1ewe7xOyLuh5dhob5314qW4WONkDUsW5qDg7iZY4k5Frzw0N5sPrHJic9aej6M
39fHqVeLSW20Vu2s0rOtcf8dyg1Q6FXL1jnNOfIoppCJRycwKNFn4mtP6MhYcDEs
rFeYEuGA+H6y+PdS+0ZmOEzMxR4Jw+KFhxBTDv19iMnoqXz1MumhhKfXvaql2kKT
XWmRq1QbqMlCoy1KREzkJBXhUvRoDLySQsveWF/M8Vg2JdNwWoHloqmaolmVw0Fb
8Qr9GnezLK3sUH5+AqRngp2L3bIP1FWiZihVgHChuH8z/yquPRbU7weoFhqviD0r
7k6OeaVycXVoXf1Wn7pANW/w4R3UvazlzkiDjmD2SbWkF7i93T9/i6ZKaOpKSonF
XVJDnuk8L3VQvkcH5r8oWnuX8OW9jMptgXuQhsnyDfRLcHZwA49xd8x8WU0l6gNd
jtasHsrn6CbGL1sQP37IxUZXgbPB1zRvuxOhlc3rMF8v3mn1T0jaBklZuv0eReRS
1G6vTzByWH296mDsZRuYDdqq7RjqfUvP1nkZXFidD0c=
`pragma protect end_protected
