// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pGgv2DrjRa2SSbs2obmwPIympmI7bOt8Gu0qGgHdKPAlItTcYL30GvQi4MP2gnz9
vJQJ4/A/Jc/3csDB1ApVihRyuV5iY2fSrCh0WZNooJFcDZM5YkLMF0bXCd+tAXua
mMUypWrwRJebX7PQOT8LOVcg6IOTD7AXSLNmb1pIgnk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5456)
I4X64A9Vq4RfZJZhkMGhcbeKgpa3WI2Xrp0bBBtXebHcy/kxPUxLLIf5KLJ7ScFH
ECCzszxz13Wyy6BI1EHPAkjc5hHCPNSUS/ZwNPhS8mkmlQl8oFYGdU0rRizpIVcH
4eE+leaewkK20TsfGmre/N0SXId+LfRgwX1MCAJwV6rl1L1JQT7mKisULQkEMnRh
IVK8HQ1FZ6/vdFDR55pzlar4gFZFBf2QZiSlFngMsAfonuv5mbv8dKgKNv4mbuO4
cee4oYc25Llr8QH/ZEa7GhNyrCYcjvlO+BFiHE1CwqvopKVTnXXJZgRaMQ68x+qz
4ouuqWwO1kG4PwYONBTpj1n1ASSTpx/IhwNxJV407b/J82ExksGwaZXrvxqr7YYN
DeWes07tsgyAN2FG41Jo1aPQVoHnHu1uomzLCk/LK/4w/tulZ4hUuTHidNaXVlnb
Z56uGp2JuY1Gx89L8093sCEXH9ZQ1qSxtAJOKiyOAfcaSCRlUXfxO71A5DxHuR79
dpblyp7fXYgz9tdoqudvfsI16bDILGLFpJNn8iSlVxhOWzhWcwDxOLGiskDCs84a
fGM3k0PRmHjzmrzM0/TdO0C717FBxeGWeTObftZIUh1I7uQ0CJqq9NTfUvfw9cb5
KIfK3FYpTbSaMr+gOrncl53mBmJnf+3L0uZM3K90WuVUSquVXTGn0uEHUIc9mg/1
VOLkACD8b4CGXJZVPlu2w+3U6Ts8eI24WJ0Ijfpz32lCM3z12mop0m5H7I4ytHnl
2vfiXX31sTwertxJB+7n/dlpBq6tol5D9fLU63BYm1r/o64bSdFHeIicYA9X3Qgr
2EnpjXq3EUlYKmOCHyeBDpY2iTTOxOqSl0imLNfCPlnVWkdAqdzUli+XN6wdczNQ
6GYDob9kDviSMBXCn5wZ5foqcxy8hU3HawaVRPfmfVxJkd5jG8XHRM8vJgOK2kiJ
IWE0Z3QglHnr3wjmAmQKu4Yyub5KI8aZYASSRSiTB+nU7SXz6tc+SBs/sIWV+SV3
VkqXPxCAVnXMucqV1khNnh0svBdZUwhFskopznK9xpEhcZWrbF5AC4Qfy1LLDTk0
+aEGJKvKBYuRFQWxEazRBhRWeHozYDEM8P6PQ+JzamQ0of7N3sWuh3EKtvG7FDVV
rXnkOhLNi1azrbSvkeCNgk4MJtvaRFdYZC4Nq1C6raqCNOzD7DGBAYAIkjXsiLnw
sAZQGQrMD78yENIxhc8Z8O6vTMeyTcpgheLMiPG87p0OxLPBiktgWenpl9JJmV2t
iqCnBxsin+vXzQ7DWwD8rLCgilL0EikWW84J6HZ/j0fuLkXwt2Sh61q0nsldoOR7
r0BSWy96KJdTTmbUrfmeYyLVEvdpwmtFYvsFfVAVl3Zm0Dy3DUi0+Chw+tRuCQVr
w0y2yQvSCE7pn89TNE1E7N3D8MVhgQtyYEWnJJJDESauKcSbQR/K/60lvPOKqz3L
ixegpvmTCFL6nn7nJ8JFmCXZydxoVgZaCbaJM2oUJmnjgjVoxJX8a8nIX4hEGOB8
GaEU1Iahu2XKWbEE0cJv8C6UAN72Csc1jNMtp+HddbLzrRGtgl77pVVriokgDztz
WtpQ7PTKmEJxu4N3mY/pcgsQaZfZO5C+ANiOKDiO5JAVt0K1LbQ8uTXnMrhZzlo9
kGippVJyRF37DYGO2LZw6xryBeS9389DG71ph2/Y5XuRjWx3/ZXRm1Y0Ykq3lHUh
8H0+sHposyFXDGqq6UWZyXg8cVelpAwcRJM6onetIsEp0LWz0X7KnppWFhdo7bnF
WYHeyF4wZEg+a3swwCOb8PvMlnVQUJee+8SR2tfQ4U7F56wg1lx1ZS7BzMdIp4mY
fMm8LQ/lHUzg86hejQlRYXvULUxqWnqkReUQjapywDp19uq28yKyUCXWR5KPkFTD
gwMfYsmnKUE5EMN7Yu4lwkyFiOUrBqO+qdXPyhtb1v0UZw1Unlr3Ra18NdStHbmJ
JMSc/hKkXPUmvuWvOxHSOcfu0oeoTRXdB7kn/mE8b+QN8fo6jEhWVucWh5uFdHVl
GnFSc8Q/0VYEdNxpjgoMP2+uCgWBLauw3hVQpKEqoRih6Zei8Jp6coPmxKLAcjaV
0ao29KHvZofREn0mhcrp1pYNXS1zlGuhDXICQjnEPJQdbPl1kL3rzIwMWwsYElwD
lsqNaIDMqnPb6SEmt8d5LCtJkHNk3AEkvVmGrhNXoV2GbrmRxLbfXEE8iRXsbHvm
LJM3tgpdP9Rm94DSvxgd55EIpk8LSa0IHw+BNDOwJPvxjatol+wNxXq/vLJFSQVi
4Yb6tikbO7YTLGaMRsqngq1qBR2FJgQKKo1W5JcxueVh9shuMrjQoIoG3wCEfUNL
GSxKuDE35de07hwOubWsxkh/uwbycIxJWAr9Frex38Xkc5Hr6t0rfLomuYyIvSyF
jEc74xjz/J5WZKLcSZrCodMkcAwyfiW/rtzyPT3uYyPxVfusamRBVJCf61jcDufG
1fEeWfKjzLUjUh4rC5ZG46iynrIZHG4BLVA4KhS70iWChpWRX28tONK5DpizVClg
JrUAjW9q1EAbuxc/NThgAKQfjwAoIo0KX9W05GCfG2k1zVSvT09o7cwureNU/Ar1
EZl7tBY7gCVzLBAOq5L2KhwTmbCoAmXSSh0OxKslyq9y8DxoGgbkXytwVkSVFGhN
uYDj7yUKq7JUP3A4/zbgjScz15ZRyvlv/f2BJQ1SblyzaPVy2jtngezIQ6BY632c
pVsAfCbhdvQ3yWSC5PNXfGtpHp3DzVpKbzFAx64qLFL24ybvj/OYhaDT98UElxlJ
kwLAcVXtmqnDu6QDhFzqyQ6cS9QHdz/HiXHv1136cq92wPQ8sZrE3wmwxiPLNrLX
2iqfMBob9P0OS/2iCP1KEf1W9NAsZJmKdqmmbelvgh2vZPM6EkWPUzg1HzRppbHI
q5lAg1ScUH6deqi3+8ZwAd7+nkzY16oogArGjqly3i9kky3NObRkDoFxJWz67VgX
Rmwat02H8oZgo82yZi95p+xn8GPScVzXCMLMVs60jIjUNdAAylpwW98JAvKOjq3i
7K095QDzhUuVhCIN1xVWy6Hh25H5uSyzMFLbGpbReqVsKdhqAQ+H3F2GeTs+2mzK
lXEKMkv4il1IChb0N0oW2dllKYn7Dwz9WHynhz3AIXiXZ0vJb3PwEFbgNjGiw2uA
LdcjeBa+8xLIZEDJ1G+ux2H9aUAM2bo/ULmjq8G0iI6Z7GndT2TvaVitVkmn7uss
xWSE4/Iwt1awpc1QnlMIkv0uo5jKoCdltUUZxgAf1EVtthJ3WbeQbmOsZ6WMx9Hj
3n8BHxLzgVHFyxGEGz88wFvkN1PPhiPVoSJ+zwi3wue8ORyVqAnuGhJ0B7KHKjaK
gwIPCYyHfY7bwbHgGhdcVqB5fjyPLeU8wN4gAxp/c7dRsrpT6vujE/r9sr/fLk+B
WvHuFM4V+rHrj+cmnYNiXis3ujvAGEpiNDRWiiZ22egAzFs1dZqZGu7ChYwkclGK
GvtCUkvHQ6L8NegXGHgStEPSDZ0Ds0Pa4gUi47z/esT/Vcin2gB+vm4mT7Ycaw3o
PCTLLERNqsHfD1y4H+UU8v8AQHBo6n/W1lv7G3uIjEHV8qfZ9oBkmhwbQS75QRmN
kQ5PeUDaiNSEG1LViwARypXmKlyQYvYPXgkDX3i+kg/Zf5D8p0ruV+cTxzOdEHZR
JvUKMRlF2VwtxKw+89L2pSz071qWiBj4ujkHPtjy0OMTmJPZWfkoqUIEKgyYmNVV
QGw6+7yDas5CgCQ24iVZ/nG6n+gxS7gntGKj3KdV+vWjI1THSFxSkJwWmRAsrcvM
Y+EPjY+ITDM2/q0kF107vphu5JpVNcGTgHhsZOKSAwKkf1wCDkFgvPGDNTGXgGNR
RK8s9S+sLiwYpKFodgAMexVtrySoc/PeEDYPn542fj98+GVsGVvUJmRRWXmt65HI
X+3fu8bSr32RVAt9QVahIWM4I/0QQJVz7zwEYUcxtXw0Rv6GhVM9rY014JesK8I6
3ngX+fxT0UhHSH3zC9s6Xdkt52XkbHtvvrlt172RlKqcCDm4POmFz3PezNXBREBx
+hq+HjEHdX4D/j6jnnViQ1gvXFtHO2pzIg22yzVjlGNlodRf7PMmsyCW/8pwMj5E
b2ztBEyCFraAokqwaj1ldsLM2MQfEXutFwqQ0u8gbICP4WqvbRXCrBTNYTbQbNwE
WYgEMoQ8IEginJWIqff/sIkQr8kMYpXzL/PV4ZdhZLmbRb7c0cme5nZYq6gG8yGu
4ROsE+egvkHdMP9JFBVTZbuTABTOTp7MEhIj2FekXuGDgDucApKo2EHcQpUyDAG8
7j2+5V3987S+LZDTXfgQL4Q+qND+61HwZT5o1eNc57PLAElXvrBtAEGrSMjFhD1E
PQsNS+tauzw0Oy+pKGbmxPht+/ZJ0vMi+3q8IDcmTLI2MuB64mH8kZ8IVu5DYkSO
u3GOkWLvgc3+QsRatI8ITONxaE6feGx7CSFVJ0XW5+0t3Da6pvZWy7tLq14jYmfI
/PbXEEabcN4dNBc6f3mwJy9LJ/1IcgHz5BBT8K7D3YWBAAVVaIsG6KDnt1T2VeU9
DNOJ8M+lwUQCnrCqEvBIkInPjEYbExqTdpmElisR4oEgjVk3FhDTpdSbQlBMoOAC
3YgZcYeocUSCejCsC29ioNSaw21mJ53FbvfYVJ0SDd1NqzheUGtJmF9Ki8/ch9hf
cQIl7ydubbFX1IMqoWfWZtKkxU0g4ZW0qybVptXkiiG7zB0SBZMgZTcNkbHI+EWU
eVggAIajSyEMO3lECniXkvTrWjpSJ3Ish2zOFbdufPUvsYxarX3riwAbUihg3XUa
1Gj5lbH56LPzIqvXy+H0RZR8B34JiNmyyJuU1apIhj9lNF9+9QweLydnh7cPKrJx
eas8ACtoNU2fluwmE5EhRRAeVtewwshI+kJZ+DOT6cqOu4dK1rZT+SUyE0lUYGib
3VHuW51F93pLqqPTyrWKGpS1AUkJc8/0TCbHNmVmRZIF0hdiTwACh00YbSozLAnO
r99MNDKxExGgyiv9x+RIsC4c5Xf2L9tdnhe3esRRr0rWqcDjI2mmdzK1rMg8lXA9
r0HnGtMOcULdCykkzhYhXFEzPwlXO4Ca2v5V7DFpxkpIJg8uhIZul8dZT6/t3qF/
xbgSpJEwW/4P7Re3Q7hQveoKPHWI0BX4t6Zl/pKs6U1mk/y51vaDCiqlgKCtW5kJ
WP9mHz0jFWgGzcpB3kf9tdOC69XSKboJpRY6/wYGjjWbvsdoTy3WjXHWQ/hwSypu
VKMGj4ZmSQULvqePOMyBqQBWRXTRQTzTReZ4mmgpsC1nVL1Hmay2M0NlsoTqVqxL
PJn5/lYwIs0SjFUX9o28vbJEv5Q0t2FFDnVh/FiEux4FteEssZ1T7gWtqWz+b9Os
dMZ5HYYaQFQm2k48hkXNFhazmYHyzwZP9UaNtQdPqwypYxHQnUtdkgCTmIam3KbR
CKPvjZ+OsIWW24OtFhYSjCGjpuBe3XruIUaJwgNSvSWUQZ1pSGCXOG6Xui6nqdea
umicixfdrJtoEJ0dsFgJbiyWATleNpgBlP+WfGRDOZuw7arld/sQAu5ar3ZNN+xV
sXKsh0fjPj0aJKQCKdkjDDxpCFSxINDGFz+T3Nmimik9obPuYrw52Qca0BAuvDpA
5khlo0jQMrfoP5Z4gURUAHV0ZrvXllj11pzj4IeIk870iTr66/h0J8nP3njLc9Me
8I10+njrD8+qg+pDfMfMgqOnrfuPnwc7yUgvBICgd77KnOiskG3EOvSqhzErGxRG
t/m6A9Pjk60RWU6RcjV3FBaPzUkeHTw7C0qsbYQSL4trrzhj+lQXfdcVgF9j53nl
2mC6O5XHFdQSFvl9fYwpxAaMGHifYmS2I00OgsBWrYUr8D4XswHeW9PbH2Mc/0mc
cAs49fs9QmPw8zPpAyNpFyfL02KY6J/gm8YBILmxLGBCkmJgslMVkrk1ueZq8aao
FjzONDOGjIwpp3vsXFRyvjJb7hyYcQqM7xKsMTB5JBfA+cBvig/9WIk2b5Rz63uJ
G4S5Iz3OtA5ioT0ka/gZzZJyYFgIvZTRev2f/pLIQ6+5U64K/FRLQjiT8L9XeuOO
k3TaRMpWBUYtKZP4nsk/j7z506kdNjh4Q7yvboZUpWFacARHMT3pxWdAz0uVIeDi
sufpahWea34UapbQr9jJjiW99Fx8xv4NMY1BB3DNdRFynNiZoee8xnbIR7Pwwfhq
D9a0UlWL3qFYqCLpT4fs/NhwsFytdHjsbJtU17ei8xVeCIKiMHMC5ahPLu/S16b2
TZZ15o1ZJ1kfIW5axfFQcp761do3TtQfWigvAs1yDfSs47orBxRixKh0XqgcaGXj
2hwYJIZKdgV/e1hAkDLUHkYZtETyTqRMEJhRtcjs4fLByoRhczKEpSMp/ivvqrK4
xCH7f4Hc8bhDPtvGlubNJh0XKZEU8G7rtyXBCxMcFa29fzC5ann6vrLIiFtcwKuM
hzXqJJPwq/FY8wx9yi1i/00Mo3dLTvCH5bar2n+OEqEGzSnLd7qhqGwPBGtgmxSB
Vu7o2NRiCi3vYBahSR9Tr8Pzzw4BiMX6JTlnPDN9XaeUuptNIcxsEeNd0dq1z6ZF
13FXSeuC3xv8LU9De3ehDwI7WwvyXaJQbvbmKtoNXKqIujhyUfI6eJGjxeqxl1XI
BHrovPcusuXT+Ms1NgOllIR1lz6tT66PNP2iuSJC3kTIVDFNlBQb0IXIRixqE2rL
wxVHge3Wacm2obkDi3jbEmSbY32lUYxhLbpLWCqILpaZw6ugzeIJaMQvzpgUwKom
KF7EdIdqv2H/4uI3Nqy66z2ncljR7UfHDwtww6lCyI2b3WQcE+V9XQc5uO4tI1G+
BXwAL2Hq7lDqsee4OGUZ/fCA5udM3S9A3Cb9+Iy1/GTP47wgAW0cHf5Dka6M4mh1
+Ccrx8VKG4sVdRixCNHpne/cDtGH0NvihzfD4MojC2vKiX9bxHQ+d/BZ9zrjXrD1
2jhKpyTdSnymD94CDrO+yxEaPjsDWly7UVCEB4U3uV4nzolbu6p5g9N84mOz2mtG
n07EswfP5C5wa8AkborZSjLGMy45Rf6zOk7jOwUfN6C2xzkXmSZqOFQE4F2esARw
REXiCPuyr5qCD81Q6Ks+N/2uMk6U99KIekOjS/AImBovFL4QgiF2nS1tGBd6IRWL
1ufK7MGah9cK1G5BcYjHiZsvH64qsjkj8qnTAWRdqj0=
`pragma protect end_protected
