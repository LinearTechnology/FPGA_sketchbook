// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lkSL3bqK0ynftw5SLP2FXyobl3RyAI+kWegj2Al7JcmJHXI8TSIzEMhNxWtHh5h/
Td6BlkSZ331Ahq8W/eou0Q/AS/UIX7gZX0V/866Mm2LddeWaRz1ckZxLhvcii8Z+
/e/MVLan89tgjsCm/SDnGA7mMPKFHhwhfdAwGVNhJkI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18112)
J7T5773EbzWrL0uZspLmiKVGtO5ypYYM4s8F+ffVealW0pezw9VHXybToH0EOnZp
7bbjWrze0Tm8vWTqjOpxAKmkCqjwFaXMDTb19MGaZdDxZ/xl3fMUxG1GrkMcL8NM
L6kgaow09GBcsxTJVeVz21ZA9DEVZApmUAWKWkglAIKic0UuNor44HAZqYoxaytJ
QM/TxMBiz+HAdpENNw/+h0cusCytFep/FzW47kLcyB3PzwbiTZxGEofwuuJM/Tak
9lcHBlBXIsbmJVtDgsIHu6gpXPiLo7v0whmEx6brJZ80s9dqXlz8E61JjP25PBAM
lyg4gGO/Z0liKSVuowktbgndwD4cTC+4s5zYVtVO9rfgWeC9cERF2jrZSpxBWHIR
O0rAznB1lGZvyPFCMRL6pQlDG1Bn9hAkwb9m6O3Cg2DJ8VBLv4Y+1NSk6pqG5Chm
X/jtFCayCESvnJidgrrO71PASEac7BvD7CoAejjL0wOcUZOgIlRFdsSD5iH1Cplb
aZFOMRtUiz9B3jcGYZ16HdIb8I3DnI0ToeomsZAMnsgWCpkozhSCQHO0ajKLe4FE
5wJKTDIzVqYBRmrufHSNM502i7mp3f2OaZ7n3bpMprv31Ou0UP6K9X5BcHy1O03t
xlbpcTxml3XpqSrIIzs667FT5CP1wlLnZofKazMV0bt0fwk+Jaa1lLAcM0/juMRI
YWGCokJTC0mpihGRt1Gc5575vL0PNdrr9fLjIFkp9T8Yr525IrY40kf5OBFAhuFb
LnzBTHB9bG+KeY+5FSO+FnXhRA89iLzsSFJfhcS1zgUCF3LDj0udTZlAcpphiVTQ
bIaih2KliP+XU3ZfnfThFDhBPn5IlekiHdbmQeWMXou+NN1BXk8uQ2enUkNonSIV
tp7z4Bibx5sum3SNtGVlj5Mv44ZV3WhIG+mwayL53mF4pZ9vumXisNglmTrH4Aj7
NxyAas/30JWh4Hrv013pP6uLIH4NMLgEjtWXh+tXTfI+hM5hS1Nq4v/8IE5IPAYF
PhriKQEcJFH0/koYj5ZeG6/IgWQKLps4DZoGX6jwi81NoXljpOhck5jRClQdPKvn
E0eP/8MgbGQKdUMIbEj2ceIUvH+gY18NnvJTUM5J2aGAv9GfOve1SQ8YEfvIZEJ0
uExtN5iEkse8BKCNSCK4chlsG/ySCFquEijXNX48s1jscw1wQJ7YSzoqy/3Snmrv
0fT6vryN8UdhFqFBGBax9Ppk6J0aCZehNy1CeIXVSH7/n+vKytJPyYKJDnllVWQa
SKlKVQO9v9Sc6EfioyYm9+E+dhRyy5JrJPgqenoRsSnEvIdc5++PD6i6xP3O4QyR
UxoFz2EMcrKkvTKaPjEisXQy7DJnjNGVSDSAtDuQrAXDfj/Zq3/NYkpiFxiI7jQ0
VoqgrY+tNU6TGD7PVwYH4/kIcm5SGgEc7lnbDL5I90G1YWQNyRcymLV45HinX31V
0gAsVbc4ObmOkAZML8GTg+DebSzBvqp8fmB/6wkLgU+d1sI7XUDiVlmn+7Rq/LNC
xiSll1kS01sZdYoashdEOPDJAAo1yGnYqjLSLublEFE6/ggT+6MGJvZe5NO8c3A8
E/LZIFe1UDxwQM0G07xQ+giNhMxIzBMGRq8q4x8//Q9ARCmyHzCtgKwtmVw+Oaqo
ksznwCmkHglNk/PYJZfyd655JeqpUG9Vt0Ep6koRnHuQI1oVTpYkINpQeKj14+eF
pdw0TsDhWYKoLpEaEUeQAZvM29W4s1c7WaIJubV4vEMb2SNBedyef2uTff6lBg+j
jiT3s9ys1noiAagQo+YE91YbmpL94t2uZG4NngxOgUD1e40OlZRsneM0fzm2/kd7
X1GCrHbaPNd/jb8QOAP4ozFtjXxDw1WGVhP2CuCJEbHlbpudfdf2ZY6QjrcPzWba
kt/o3wGV9exeIb57n1G+Uj/hTbWkYWUHlG8Ha0OUBEVUDFj/5agrrU7ok3IKDdEn
mxgTVPzf/M9b6OgnP7w/zin6xqXxwsMDTRtLNc/yN3+gB+YoWzka3fjhNNe7JeoV
5rDJBt0zjYORhoFiZirSBV+Qnw6DUuJ4t4ladvfzUd11bi4oiObD36J4t8gi2Zqe
qxt1z80KVYEV+m6jlnunKdOnoB7mS9umBM+srd4bQXv0EIbMj8s2FCtguBTbS9iq
K1El2pSuy7udstOG3xNiXuTImxSv+2vXhMhQbNT0ZJ9vEqMtlEvOFOkaUHE1aj6k
A1wifa9WtvImmDCA/LmfTRc3kBOJ2PDMmmTeYRAx01Hu0bNg9AriqJBO5dynEgLJ
cDw6zF/id1SvG9ldjHdZQzQ21g8kOQhYP2i3FR9JZxMUdyod3YLncgXxmhnuNrON
cjtrKgiVk9VXT9yT3PUo+GMMM/RghwDa4i9vnmxclYIJ9yfvrRIw/6Jzbzp/zuGK
CpSHKcOYja0ZsMG0JNB0tYha9BOl30n5l7/27BlGr2HQ6xxzrPmfWI6H4ZXILbR0
KKvYrZvNM1ReJss9vS4Z7J9irvN9GJ0YGsonfDet6V1IC3TIGjTby4WySpe8p8VB
bhHNbVBTR4YeyGPhazD0jixoMxP1PkO85qkai3+12im4X+Ng2DkcBjUevCIgl4aa
4nP7ePPONevLBwQYvEdrn5bCkfXM+sz+8OKN0A/1zoQL6sqFUsG/se1PoThFURYx
JzeRgYwgDKPGcO27VJ0QuhBJFs6kJfUJLpmyuXUM3m8bKwmKf+v4ZhVvqom2yxCE
y9Eic5P78MH85AhoYV21ekQ8jhmydacFinLeYt2P4x4wYcc6ikDrxQFe9oib4Hfg
seOhGpj5V5024t75L2heQUQ0AFLTKUXGhV54xxRJddhQHnTrtV1owarxNhHVH0yw
e7g4DsSZ56RjxgvbFbBvpY9xLeEw2SW0/xabwkBvqOM6wakNKn+nYKNVXittUIb0
jGnQwDsoLbBATTjwj8VaFl5gpOofYnkXMgFza3sqll3hQ6hKyxs0qyI0E8l/3p8F
KwDaNSCHFyGYBExMuggeIP7juPbSdQTNUqD2Of4jyN+0Z/yGve9owyryjS7Y12gI
TCHUE+71uLjbkiHoZr5J5RTvU1ZSTFBrrsj3YL3U9YBj8IEtvGcPcq48KJH+X8Ev
tbMK+hOdJuOkqUBe5/3qtsRHPnQkBbdJU9/sERmKtTbwK6METf6rLkbM7pZ6vcLb
gbGODiTsMKA6piVJZLxoWa+NRgHVLuwGsAC15LUkWTkY+UEbqOZ5ohQqVfoxIEkz
dhSlh38fcBLiAIr1WfQ30ybXZF6orKMS5fAX3nyoerVYvJCkt8deaaqIHRMhd1O+
pS8lTfkJYX01h2NnVax6HyLIGVzCLyoCDU+WG/rC9qgQbpsrlLxF59xWd9V2zldg
eIbLBW4lDk03uLyhqWwqV70MjG9bseDCoRWWD54rinFVjAVt2X25CN4ehI4RUPsz
fJMLPM8Lb69DzDh/VKBJkDKuzLx7SuNzCTTnt1YuHa4ngfTkb6CR2mN34a2Wi5ZX
0uPjlpBKbhqft3wbawCpX/tx5zHywp2ozn5vocA/czQgwI6FIoJMNuAMhMwcEQn9
bL+q8Ib1dEb8nxvwmhTK8gSJx+DcfNOC0sN6BCdMbKCi9fjt2LBNrXELqjQ9jOKC
A8lE4DQrPEP5taT8A/EVFzI+eNublhcDMPkT3AZdzIixm4rNSU/+LTfME8dJ9snP
vCl82HkDp5bfrwVN+CaW6XjXOOPRh1HfDdpYeA/DXjwG+ueeKs4d6ZrcfFQVqQ4Y
6FdOVHQtAOaSxhE4PApyfnTlgbj8iUO6qBLCR/6HcoESjrM29ykvq4fO1O46oWPn
8BchqlKg8XgRscdcOKcdHrSBKUxMY+g5dz9IpHJS3W0Dc02GxgwhfaCorzj76z1H
1Fe0DHr0LTbyFcGmG+IuHm/VnvVOXt/kMqThBQnTYUoLqHqccVnkVnvca0bDWQay
WMTYIO+U15xgcH/+u3iKKFuoblhEqEfrLK/V3+xY3MStZ1mxoRPJJWdtGrRY7jkx
fVPxv0PknZ9RYyx+HyXjzTrW0iX5FD6q7wNPtyNZZFQUd9l3q1uAWMirywz8LzBN
6mJp/+NoCn34A9QsGv+fiP3fxI9GQGOT3+yAX2FX35ouSHMe+6aCXyA/psU+6ILR
7hnt7erjd1bkJ5l+WAsWLP6nT7k3U51mIZqfhzw57wRwR6lXDrpyATYIsCLsBm1L
K5ugnM3Du/u9+E6NSOQrYkAVIfYOwrMcg6q+wRRiCMaH+gvKQaZ8fsRQ73Cik+SA
iM6JwW5jGy6THk00Qt4mpLDi5hxS0Aq7u5TKaoingV1eNRXRIBMPkrPemJsHsKkI
RAO1AvUePYKft+TtzrbX62iNCEuy1l/GM4Dk0FDpYNg1H8qdthQeEQ9OPAf7IGM1
2ofS3DhH/93OA5sVya+cS4l9XPCTO3MOqkYht9TvPPEsPJvbKbvu+f470JL9pihV
qiJUyhYh5SMIc9X8OxmBv5DeeTNCgqv/8/pQXcsYxFHkTHYYber3/mhyWNb1+oVT
YqyL85xCvtC5X1Y9dZF2PKFzr5ApJ5q1IOb68YoXMxR7A8iWERfUALMBZjefixo2
gSBphUxUFVn3V2xG/7jBvt2WYubT8fvFyEiC4BJTLOixeFhwxQXwaZWzSD0zE6PK
IiFQWpwSQaiTvXWH3FKkNFy8K5cCX/b+i/hYn9Zsg2CNBIWbsISPEbxn+RrsgyhC
ZX01HiPE2hwEHkbOqXtaDIqPpk8IMTTsBLy3HSf/zBAsOk8ZzLUDVz4m1HgxG3G5
F5NOfrwfz5hYEIK+jlrUaO+xLaNuInqOCZ76bViNVoj1IfBkO/3TObFI9nh8m1Cy
V6cxBDgNZ9aZPnT6NlUo/+gVZDPG26cFWryQ9TaPEcZfFtBok0Oh/WoIihMSbK5K
vYeFn4hoeWXJ/aIsY8GXKOJD0qPLT1Y9zEG1A4uYG+QicH8UZmaoXAA4j8507k3W
e+PNYlc14EclEnOxszm1PXdElzQ44zZxQ7/hx4rrt+oggFpPwDBTJiXLX9aSa10c
FEd5sHtvRzmmjixVbPCzjv3U3qIoOsMxuRGCrrDLG/I/jFbvtZVijC0orart/Y5C
seWgxFBR6AKvqu/lqluEbqcSRjLoglkE6kTzmb5JZCu0Y5kzQFNwB3fGrLj4s2TW
Zuw4r0K9fEB3oldhgV0fheZcmNuDXItk8XKlFrIYhotmOlrUzfwwck49ouP535Ae
V2hlAwKokSfLDRN/YRsrA+8Nnwq5mn4JF+a6u2686Z1rhl7MSMBwaa8pXN+EwhJx
et1Rkr+nUBDMBBvhggZ/KCp5eDEfacLV6ZDE0d0Y5hrtVkNqRHmjAzi7VE6iQ1zD
oGRTSPxgz+LTOsauGf7eCLL0EsyPvw/nqMxa9+IOR0q0junVCY2l+l1xsrOYN6Es
iSiSq259LUvvR6bHeEAK+4v6uRri80kRYLkGoo4Ow9zsHBP6bKC41mCA7Ye7qgYx
ryuK3FpOe65tLF1JSu7KnWBrhUjq5KhDoLNx/EpPCEcFNqOLI4YTdog7Euj07Q5f
H8IIOdieeHL4kdWNELwgNwz5Qma14x+944a2FdrDeJbkDstFGc/0exltdxb4zWr1
28GZNIN9vOPcggwLw4ljiyb2IvYNz2ql2Oqv5DlEvPD6UfLLU+h8FzUO86j+R6b6
zwRAoRqYauCvydhg2bxMCkKRRduGENi1v7jY553yxkzFrNWrw8jYdcujdRVtnt5y
V1fvxXllYECRUtn/zAWSTMXSp+8OawyZS+stLiqJImNRzcYMf9fKocUfQLiAVuJs
BzfdbTxxgr9Oyu2ee+E5nsMygOmfRuqgnkcK8ISbd9NOB310Q3aoC1zZg4CBBFhr
CsozvqnscBKrrZLQQb9bY31tVPqqTFOt3kKDBE55G2mVjD7zvF4d7eqRuXI3ZB0b
ecFjtZUwath4gA4jNjaV+gk1v7S7VJSOeZ3VhC7Z6FqVNnGEn2sk88HyzsTSh4T7
PGxTSFiZwJBeC52jdUCYn6iUGqO07E9MMO6oF2Io/Jn8gziTr73bIxrJwWcxFF5I
GIhKcQHnTFfPOkceqbVSgBeG/TgaIc0Z4SLhvheByXqdWPnBGGPk95nlhrHLGh6G
Um5NIc77aKl234U6jJsylKnvjCGD14gVQLB4pwCN7VhLZmwBxoA+DJOpEm3KZWyR
QqOdhMOqL/HHBJbAElLxZLqlwxPtOuFZJrJq1B369pQ2dPLzFd/8sIk7e4LgoQS6
oDUTtMnQXCI64Da2UtQeHJ9xf5NpGZ7cAKu1oD3RtRGWe66DdeVS1QMJ3PTYjc2i
3cFxcoRG1yNZY4i0ZCvO9T2SoYBYjG404Ps1Xf/McvdkGLXc/4ElAqRgY+7XMhP3
HePSUulTjA5Yoo1PEq8OiProqeBwXX2lxkggz3GmszmjcGC9PpE5VR8M/pwp2nhJ
H74XEZ8KkPRQ8iZIoKpukl1SZNAFHtIw2BBr1RXojVXmNjBySgaPf1TpIXiFXwpp
CW0R0dnEvxYQm2DWVRBA7uApYdijdgSCc3n/eiSN+OxPylQCCmZiGhXy32ht++lb
0JD2tOb8LSnXWFdQ4vijPlFk14FgzOXvlVEBcAt1QeyiDqf9sjsesMTH0i44MTuv
5lvt4//oVHJCef8MvD+9ol7E6qzvz2l5woga2rN81/4P1Ew0JvOSv1Yq20rNgN58
MFnLlJOQ9GVurD9rxFtzS3eBOoaXZ2cdLyi+kUcjzRF/924hR7IxTNwWCIPRAgh2
mK+LJIuSGMLOx75PtjtYwszx/Onh7zhXcEFWmELtt7MS+pYikxM2wZ5awrNfSIUj
VM24mCqA8oWdLORAMIAQkN5NdJKbU23PAU3U0XHx+kxR3mds+qBYwW17vtvSc/3W
vsAVQztAY/Ar+3c0jAdKsNFsmv61dokDPpXgQ2Qz0fj5YU1dAFEq0xsuoQjdhWHK
QbOCOj89+U/GGpjWAgtwW3kqYt6aY8lkOW2uN0NvR+rhiRU1dqgH9gdbz0eREJYd
Eajb9lP1jecHx4k6o0SpsJUaYEEg/tFmt02oF/ra7GQglYWt8vBRistLFi1KDVwN
8w+g+LSu3YmVGzRNdzAbatA6kTylXlgAlJoU9qliAM8wOHC5MUOtggIt8/ee8k1k
g/4nirAPuyRD6ijtTXipyhnG8DhZ25au2H7PFtgJaSDAhkRFqC3KKFe0D8u3bWq4
1m0pHb6BiGJGDpuO9RPEZjZYnBzmE6f7oPyLWYZuQdxtKlKTWO/ckpC1SGQ+vuEL
gkHWhyF9N+pJhJ2JFNMiy7mc44p+Nj+YqnR42fmIAZN+kO5SzsFbfriOH3rF8Y7G
F6SrkEk4nuWIAW2QwgmAU/rCu+OWDkSC+n5efkiwTS7qOzDvJc01gK5dfYOOGmk8
2Dc/QrCEUE7vQqEsQxvaDkrUAyGXliHf0RFARf7d/gOdPmuk3N3YgljbGon24Ws5
OPJHzGdFk6nZ/0LkAmY6NlSgvldPQN0KFAG8VASavVLeQkv1WZJFq/cLXtD/giZQ
6euO0ag4v3pQH9btXZ3kQYKNIgPYCTe/Mggvlmezhtryv+EWniWA/QSgHgm2CveL
dRThwFwfp0Ku5R9CxjqeKbh5QrYpctC/cQsDhQQ2FL7qYs61l5mhckMoowNn/zly
c8nRlczFNKFcOKtiQfPK604zI4qnmVzGDeoRGXswITP9MZGE2VqMDkGLG0DUYirm
o6YfLBqEvozssaRg/yFAhF0R9aVwqQCNRCo4l+n+z+VkTkLw8HLAkzd14ybXAaFM
DrnEoUQSa4i0iEc769ct4Olyv/ZtFueJ2AwPaQGAZMvfL94BTVWbon7B8ZO+jzCt
fUXphlnSJXeizGdpmOb7SX4JmibdDv0+LpYbi5Gwui0Js8iKNQfaRK0QUadxFjVj
6QHOrx/oFffVMRDxPguenmQRE20amkkVR0fcYWi7wNVfW3pzk6n4AmT+omDtqMYT
PdRHUgfZNr/4S5CNUHvRhKhfH1M8b63W5qnmGj9BVeDumKHvUBYqXLVk2etiOmsq
KYSbKYV1yRu8fDfa2/wU4APCmFL6C4WWz6ie6ecEJeOBvaBmECN/Q2CwKuUKk+f8
9gAYKQu79TfL1zXJlazmiqZZyVFpr+xLbECw3ZdSqkYFHPs0grh6cV9Z+RqYa85r
y6k8FwnARvEuAfmxUVOQxodcB8NEcNj+xMg/zGLREU+0NH4H4jW8QTFPAe0eJnbM
tBDSRXUEyP8CUDkhbpgMoDrwygOIg5Bgf5wwaOZFuz4Q+UalaCpR+2mBWNVqrZmU
OZhjtWSpjPzE5Q5oP924a78G6OQQJ7iM9qN5ixKy7HmyjAk7FgwPwePWHxc9qigV
Tr22VgzRNeIQwjqL0/Xs7M5irEFhaRQI1ykgakvThVO/KgbC4kF2CLPYMTl9HXpN
wjnsG5sAhpKqj6d+oGERv+M1KQ9qAjfdoHhtCv7o7OUz8gqaD69Qhgm5aAfUROQ0
6DL0xUuUXy8NZ2PMZme8FHK4zYC7NOxcCEKPVqOGgJKnsLJVFWpaJmtdZ4o+UqKM
o6FAeOzCPaBVKqunqdaiNUJZqRnHFtzaAV6wgRrbne6Wh+j5Zj+U8OPZS1UpEpN6
R+MnwhWYs/b2HX874hlk7T3zXSBGCUm5e62lAgTeLH/Q1zXU/F0uLG4LURGWEH7v
OmkTzL2iZ1pIA+9neCXugp5JUj3+wT3fFbzktnFsrtOQphyD52vOd51DRmvhhjjW
GOSbgNFC8aJzwm4G7b2Gx1NmpahIpnmgCjpl/UxNd4hvYQ1lrTdj+vyQpoiAhWbw
oyooxvg731Yqm+6+Q05C6BT0IL3Q/sEz68VS9BdmuNrIPQQNuvmBu+pPCNuZ9fgR
q5fRgp14DdmwaK665zVI6B4tgp2BiS8/HV4B97lFofRcXyoZSjjJhpB5x2wvOmra
GVLHaR2CR7vzy6IifbaPzM0Cz6ZXu07HIsu2JpsOk41AYVAYqS695H7b7Eqv5aru
mBKjoJXTiCFedjVC08Xof0R5uztzCjorchgNoKxO4Uqq0af/i4+pUnXwrObv7jNN
N/YzvtZJl+6ibipifW6H/AX4+I75dwz0N/+dP3EXr+c7xVMLMnY/Kh+9ZQpmN/RJ
Pw+wB8w1SCUBTPuLj5tZBWiSDZGJwCkktnomLNaR4xCQAo0I3yWh1gCWv0xfTWxV
Io8CxI5vB80BiyS9Bc/Nf8f0IrQSy8BmlLxazXaMRlQG6ePNU4WMc2mbiOeJmmQp
SpyenvXnTFyK6ibjuMSZzgg10our0qCGnVpbM5IhpSUBgjzh6JCDAVK1oN96nYt/
f1HuaGocThmp4dH93qad1GgHleondosvihjqHjYPbbaEeUQEBhjZ0bCn6SAVFwFl
VMYLDNoB3OjrbsVJP01JmOHsSjyG3YQ5T0XfJpaASJcOi/DKOkxp4kgE/uWA8kwQ
SwfMgnolyrwZgVzRwS/sZwozcRv1iZqLSjBD5P/MO36d9bds8HAYjp7WuylbQfaj
vCD63sDdksXWirlQZyMf4xnvc93hne3cPL371qmeLpOR6SwE3S5asYpnr0i/UYDa
Eo8Ihitnz+C305Km94g5eJWHnbfksg0KRyMje6xdT8anfmGdrHJPlyQBUKeS4tVy
yhPhnvFcv5FtQjJ+/lqO2OIuIZm9o1gOuGWggwe2sXtW2k7E5umxe9NGZn6tObED
aVWjvo/3BaJkuVgmWDef8L0xoqZF4Mhu1On4tNFVj68cMzF0By+GJPw5S+LaDFq4
p1J/DC83IA2wZG4bmiSHk7ZCXEWeKpNieY70plpJFdc2KRsni3BViZM54s8sQQmy
8mGbZarValfPM29ndr4B+IXonJBEP0YHWH1XJGEu1QicM505guof8MUkPFhYm6J3
b6F6WKpeD6G1f3mUD1lnEtijq/6Yym9x972EUiZvVVptoLEpsJ4gQKysPUoCyCbR
/oZWPw0zBLLBeHJH5q7OVHLFcikNOgVVmX1Z24X7GcJQgGV3jkNOCxJ/icLti8SW
1LkUrfG/zdCq7P2ZqNBzo244FU5+vzKhdhdOn52cDPLik5sG6qZQE2KBfutz53mK
QXrpqyXRIJwjbvk2ghNOZoZQhC4fIVk14qIkijPxOgu40oEjVJqc8Iglu74ywAGh
/XJtI6WWGAIPWQYj8u/0PNMbb9xUvDjRxy4BiCenMsZxduGq8iYWYN4vmY7CsqQM
VjO7rzZulpQ8iZt4ZD3FwAwNYTuCIiYruHETjaNoAb/XaoxUm+v7gKpOkbClz+dY
Ki+UycAnH0ZQQ/gF3ECrgiqIVG1Vahd3WSZICYj2M3vTS3XXx2Zz5pXlo36qIq55
WzfXGRzPUC/hzj9q+IQ30yeA1K5HkeVspujg0XLuPR7+i7bCtsEBbMpLhli7YV/a
5YeEqMPyO2TEHXz94RGz2SjLDQerQUFct1Nd0j24RZtxwRfphMWCH29qxo+71mwL
Ik7ZlGlYORkZc17ZRkbWgFfML8kmnBehUpxj8kqCSPVfh+fXtqTsqjKwcczCOaOt
PGd0FK4SHUDj2/IN8FvAdoP7HrynZxIQaQnPRqPx7mtxhxphw/51bVYJIQzSFqRn
WbB/XU+/+YNwckkufdCBIhcLteA6xAgchiNastU+k7jDZjJq+BqOPAvbUneRDKeo
HjBfYiX/vXksOqfKEkjpD88G+32I8dVfOuIID5oMI0jBAM0YrQqWVQfnCCX1U+nP
RHf3HhKSbh/3e7wPvcu+406MqQq/YzcXmHIILcKkihmg0AsAynf98YylPR+9It22
t4hNTXeBEeAvXhJHcLtrCIy2d3Q8tnc0s9QeSN73k6t1zJehaEVcRtHlrKVJB1vQ
PR7N5a11zzOjdaUtS3yLjILlfwD/yQgauHLUiVHedmVjvi77pccNf+gcU5wJRMSZ
yMRXgmlObQsse+esHKZrtmqS6h9gVVn5owPCCmjGgNHFqEjcoaD3WDbUwPIWW/3R
qNa8XFdiQYcl1tuFEZk8WYJ4ku8dgDk10fsWdg3ocp7oR2WU+tgCq4ffMjZj+GQd
YB1h/aHA3gpb8/RVLHQsN04o0mFFLz3l2/WMs63ZO2EQwCNI9BVqzV1dGSnjtk1t
+aPBkYEY35SWupmaTXCUK35fe1aMSB4jJXpn9ssPzxGxUa9iBZJnRHqR4tKSYuds
etloEe3uh6rxu+ctUg+05RSo2NUI73m2eXhlClLmNevPY9GdG8DOb5nbjUWKd/To
rhChWUCl771FbnaJYE7/htrj2zalfZE8SbMx8Dz9f3XudYIW4Hgo+h+9OnymxZ8C
Drj2FmklvlFHuP6l9rDuk0VZ5FpQ8e3auN7J4gcS1STnI3jOOEAUTSalIlyp1W2M
GONlwoA4qgkDd1hMG7ig1zTWLDdDopInF7rJ5AWVXYEtNWlgOSwBaj0TCAaWIZul
oEkaZs8NAId7xKYfp1EiwtJzXcR6KJ1p5Z5vt+tyzpNdcJIC+s5jlhVpHLIUZ0jw
8xLm+65ZeCO+KRPuxADr/ut1oWf29VT5Q0h5bpUZ4JnkdvjI+nXXqiDjJezXCdyp
oYgdjuntN67tsnIsC02bQ65GkPO1BMcyvLw0ZNeFi4OLDqFQoxTmqlJruWPNJGbC
eFW3TMAc65TK73J8B3s2Wn12JZx7M4AseLjNyvgZDhFd+lHLZwh/+BPyXL9KTczI
xMRXQD4rVPxS8ypAuwapxmwJEJvkeH7D3MkvZSyKs4x2nhmnjSDiLKs4/4PHwRWe
3S+iKKGGSos9yeATYUheZTRT8QZFlNV3U16nTRjjjlk0XhBQAOwIVquj0Z3c9h82
1TUsFiak6aAzSq+b80BPJasLiug/n3EI+7+9V/dWhkoQnsP2A0u4Ia5jpe6xEJF4
bg+qcYTdF0CuPNswz9i7dPNGnlAQ/ZL0Hf1/c6kfKHd5duKhqYHehTgQLodrYZxs
0LPkXD9x3WLoe6fRZz07humlSXf8H0SMCl8JdQfgy22SqCsXgZccVh/iXZ1+9FDL
T3Uqig5M6Vp3C6XRsM57tNJQJJF+VMchJlEYNHXhhKjJybn7h1+Zf1F2DsYR2f7a
1KqY9XE4P09zM+rFX7UR/AEW22ALNoabivzPqR/BMBCuL+FVHROq9TK8hoQEXOzx
2Kc9xrrgNA2X7WvYjNh3PdSN8kKvqjA7ZApVooQtNSmH7tCYhBIzqRrUzZDWOuKH
X4t0BGSpiKsPIcNhi+VixernG6cta+PK4jp2Q0wTCb1BBXiELU4XGlow0Rznu9Gf
9hpml5sQkqLo2npDM8G4Q7yvxURq13udtjyCxK6SEbzaVXViBukmunDG8ZAQDuVh
g37o/piFVJqgIP7ab3yolPp2GhQdonc/ZKfj+DFLuZuCTtAYw1+NdkClv6XVuVT/
7XT1yRV8sLtsDKXhZkWuQdhiF3pVDUH4IEQTAKdlCXfK91WBTqcvSn4vocWNr64+
0sSYqU7nzEH3/dPm22Fzs72DxMnTyTTti7OO7ZF3JR3IyFjE7zFfIkWUuDyexD9U
Pi8h3e6gLX5gFsaGxPVMQ7xP0wTp596VeYtJJxWNCE34yRtfIw7MXX8se02eSQfE
uAw7CXksBnBsdxL2NP09rDBm2xHE8/aMiVc5gBY2AhmDJZKA64diDOBqEWgwDwvd
S9ndGEpDQRJ9yIuKXck0I33Ccj9nNY5EIu7GyM2fdq/wpMVbZfwAbVgCH1yl+z6q
AZyfqYyNz7T0rwvSsX1jvluFafTxgkK5RxQXZ8EyG/JQNOgLviBb1WMKd8mjVB4Q
+nuEgk7vVeLoP0ak0UM/eeVQWcwpbvJ8yaBobQrS4URm2O0Z+RYTR+B8lQeniK59
rwjGLDryRLdSnzI/viJ/zjJAg01ZnTFCcutStVEvjSZrdbpIZfeNHQzN4hEO+SKm
kxSNeHCNM+M/03W1Go671VWAdiNJ6SZje9YbeEE09HRlRFNXexmwJwGeVQTuSaHi
gZtj0jE/lndaT9scfrxpnhE7cZtLoAgdKV3FL/TnfnAQo3Wzf72MVabUzaxQNlRy
0X8TP1pHrS8v284PAW24DDY36gQZ57RmKQnCCGD314jDcQ5N9hobF+0EhtC83FRC
9UIgbYYLBPDlgv+6vLHMX42PvBQwTmDJzZ47YjMqIYE4eTs14bSTcVsaChU91ih5
BQjrstXijp0+uzQ90M7fYr8ESFXpJKktoBjGXij2QPd0c8x5cYbMfysKWt5M80R5
97RgshxD8rUkZvL2NLyACIGTPEAHGrCeDCnHSk+eDGposcNj+QFAJTg8LftkEVYi
KLnWiiI4wddM2iaWHx5Zx/RRJI6d1Cx1weIm/tp9miAsapPb+4m46WhStPPXAl3N
sr0Rufq4RAfW+fYNotA9X3wrW8kOmOMM3AMJuiOSpVbcWdBUQWcfm2/a62P/31qG
7mqhBc3g9VX2EAuNSRPvw0BkmqNOgJl6lxo9AbxjRieAa39t7S5mVRyzDRUi0+Iy
4ylaxY/667whfV1D525b5Ko4BxNdYcZRdKtGBxKwxalG3Hp/wpYaeoMrpafjbsoU
RyoEYxF0DShqLVc87FolUCQDaZrfYU+W6igPGCW+3/xf5m5TVksBaSJ567nJFSWF
UFVSwz7nWjbCvz9sgFWv0ZsLaxsfHZvFEAh8JbBTvSL9Ni6kjIX9iKe0cOeWQi1o
sU1zflY2PDOmF7wMCgjWXsMi/D7TeQJdU3q3BsOumBVQN59DY9WGFf6m9h8SUNjU
KGyDxexmafd6MlNXNDagVUtHvc0aATtvNrR/6No52/tcQH8jle61O3XR6PyDUhvL
wl2Te1P18CU69ix6QEJG0CLNQbWy9x6aNdJ3I+3Z9eHR9mvAouifdz+a+1h9DSWi
11/OHshl0UmsZrYhQkT1css8RlQYjtDWV7OZbe6J+FC3uVE/tLeo6zvs28i1b42n
RroWeRUeERDkS4muT6GWKHp0lsAt3KoyRN6tfrxZ4YD0QJnTiqs9V/xeR62sPoxE
cGcOiIA2dPd0VJf/UdLubefus4a+2Z2Tc8ExgfE4smUjHNU/VQjbN2Ckmwqit0K4
NKU4WULRVJp6IvjLPtbhB/Wm6iZFewTArKw59tt0fHcFExqKCt+6RCqQCi9yWrkp
tUk7hmaCf1ZyNvPDgwqe0TnoI8h6b0Fypp3RqPwdaf/WF8mnxyHXyLOaT0hbvKoU
XiZyzNIYnDiPKf1axU/a5ZUVFg0AQJ1n0BebN8LqSCnP7+t9X59rlGK86Rpnnzze
oSlm6FQTd/FPaA4Ik1Aesmgnc+9R4NCVpVgOlXbrOGwcE0f/8N+81AyTmGOs90Pl
9CHbdl3RYlx56Sn+3/PYeVhnBJYGci1IcV838Rwhy8HkyAPKsk6aEw/9Te3/uteF
02KDr+sMIKGqYsTRN5/z8PiyharvGOANCrL9FYNfwiiQOZbwTjY+3+fbqODbErri
H/pX709y7Zf2sFjsIgfoLvbnOXiBqpdW00oDX4x1b4b2jnSRf0eDtbCPKZUuJaYb
LASqyZyZjfLwyePeXFtVFVTechk2gAYIEPZ+Ji1hX62hRY0gN2y8076YBRqLcBPK
vpr/QbIDxq1Ta3srlJobKBzGivTdWGBmKY441X1HxecRA91dAbCCrZsg5R7SKziG
m7sAehFINYVxz1T+yMSsMtOiZmZCJctqpwM2OBAzn07KtbmL9pGnHglhKdR/oGWw
zWdxRxN+EepNEmvEwiyIEtvX47ksS5LeS8h6QvehVUt8/9RpgYzHkilaBbdwbE/t
mrGNRFUS4iEj6y+VQBpNpz4j1rEk0GkGKUD8KOv15O8FP8AMQ5ZyTll/uEeIXjBf
gOPJz8B74rTmBfPDUIf7Z7MKP2tQfWRa8ZXV3hWpYbs7d6jAk7kOH3s7+PlDpkwu
mnoEjXtc2bDfkkXr2KWa+oJNMYnF7SjDtQkLTOWLRMd3aL/4i9+TakhwntlbnOGQ
4TS3xY6x3FUP+x9O4uNrGA3x8oKRnd8konJbNm8u+zMU5qjV5T2RIUFgut3fkL+C
9SLBPIEqB1auibISa0Qnq9ZIbWMJpTbJ72o9YG/BXCvZZcUERFGWjbSkCip8KfxX
wvf4ne98qHprD1CJCcsvev9mgWpUJzNqszd9Nq4bI9oS40p1BivF/vsmBEBlDaHo
rtBrCZ0ohvj1aeA7AQSN/aANGhHlZ3vcmZmQnwhnISqkGaNK+2j6I12fosz5PwZ2
QsupnW2rgZXmPEizGFcDO1girg4jO8WGmYSTKVrSnTlKbaoXUtPLKC/bZJGHgFAN
EseCakmkNutsjARrD4Cl7OuKtq8ukbvtYduhivdYHG/cCNyIFrEx+M5f5Gt/fExX
6HWnhS0+If7TCMw+sspqhlbp1Fft3ju7Xas5gQ2QLnI/uoUtXWUO3ABf7lmGCLkT
ninc2ZmVCMLRBtCLI9LwTiKy0QmfNlAMJVXlLkZZhYRmdcsjY0QdpfzSK5XSEj7j
LVwMaLCfQVfn8VtwOMhkZdjcShd1TG84G2QEgnvfe3liAyAEFwVxLg/tRsmIENJv
3jEFYpMaKEDnZAKh1d6RhVBRVjCEIlBVG1nhRp7sJxX2Yq0cCOWUKNNFfJ2RsYPj
7nrorIjCAqCSOI9Bhn0o6rkL9yiu8PemG3NWoxxbrSyORgvZo+9Vp2s/RFONNaCr
1E1yBcPBviaEVwx73jCa5iw68HLkUJPRaHyM/iPZaGXAn9fK0a8gDpXFFhI9oDNR
QIqODykXxOcCjB77LeSHZrgEEhd5QZ0MowOfzVnLY4lfgnwqiuFCd4c2w9SeA2yz
I4rGVIMzSN/xsCKr8ullAN3O41WGEma+4Dr5RCTC6e0Rfi9PwIJ9IjeSsqbQdLqu
m9NVA49Tcuy3tXNRGW8nnizXiZvQFEGBPvnaL3/X7BoMlrGyFU2mpnqAUt/jP9cK
aNaxLu9mrC+j/dpT/i15QMELmRykZw3pqoG8HEp+TQJOV3P4MIDJ55MyWlVNirr5
/zhhFOg4O1rNe47EhqvhO3dFaiuQf0fjadT68VeZLGFayl8LvSo/C28b/mt4CKwL
0vpWDbSNKN3i7ekyvKg9zp+o3jX2bWoIyYy+xn1QthA5mD2FEBSNv21bgAduok5S
Tz6gGe0MJV9UKJRZDX6EhRccl/gr+yUw1C+32nNeqQQRUtj45Ekjp6qEdZ6zI99Y
OVZHN7E+9jVtwNmDbQGYKyp4RLGYzHcUhk0I16L/19gZ/6rst2bRz67FWhkZhEeX
lVQ4tyiClXxK8Aqmq9Ukubh9xqZOgZgVwyntmSGlp9TN3RRjbxIxgS816Fj16h/p
67oB83+BF/ySuh2OehLtCLCH/0EdBV4XiRx2s5Tt4wTjnjtxvPrymZgB7cp/7Js6
UPVL8/k5fIKO4heYBZ5M6csj3Jdr7lKicHgWc0zDnijZAZVzMQIqaRtuAGPQ6sq+
i4NxX6nFizd5+/hPjkDiVPvxVPLIOo/yqRCSXguFilmIpMhPQtzeLFh8K7H9EwAd
lxoxLOh7u+NbphYO3FhRyjIc+ZV1VEsscQS6aDXW3fUhm6+Y6Mtpb0snWT9xmnLc
yPyaxFirJq1IIlaVg5XStfnfjO2Mv03+MFXDmQS9aburFWtyndO8lw9O5t6cssaM
s3BNcvKiVipKOMqNHklX6SPnk4ItYM/L/bit1wH02039c+72pXPcE2OalMdIce4y
cYa56/wWWVz4m/SR82eizJhoRZdKrgPY0Fwe7zKOfAgfGRvaSV9HBLiT8wKQRpRZ
9OjZVzq1qM/w8iBcT7JYrtITf35me7EoclEUWyRHGtdrBWTznIt08in2owpB4jGu
Jt9KHP6cOjU/sllx38psrQMvz4D0rZHFvpX4lAh7edkx7VdugoF/frQEwXxpAVZt
35UG9NpXZLa3s4HC8/MQDmOclbROIe1ydV2HMLalBSN9fae42zh33XSR0liAiIyz
o1WxXaxCMpT10JnZmbQGTnapMq5mDh+A0LOy/FK/8A2RtIN1bxyj/u89wHxc2dRK
e1rx9byOgO5infUuxafFZfJ1ta3a7OJXiR5MZzI9nHhdWy2MUwiTtABegnDpKZsA
/P4vnd0Lcl2lMRYnnKDh+uVYyRKjNRoaxvNOW0wa6Ul0h2K7EEQCn1IE96MksTIi
kbLFxP9xySV2aJyHFgzL3aqcjyAFJfhJ6FMayD2qNy5Tm5tc2EEzoAMYjMqQsmah
wS3b8HMKv6HouB0STKplw/4TJpPxojp7kQEuWSbPu8yA1e3dEWzZScXaUKHxC5KD
5fbgD9h+yrcl6X2NmS75B9IVpq3J3wHlii0Wzc97vjYQAThgaksZQ3ll/5QoNroK
qhvMLZphhCwiQXCvxxx+4zr6xP/eaFcBmXexDqKEzDcet771Zp91y68Dz7p/6R/A
072MCFTedQxjrGc7USZfV4IfmuRsrM7nggO71xVLGJlXCvWrMBxRz55qMgNXUXL3
GavshTsFf+gcfUoDcYpA2Bh0Du9pfkbJPulI+XA2UQKla4xcoABOJKoEHcVlzI1z
eAnci0uObJDZxm5opuwndaW+nLt1dESmVsrkn1OA2A7LyASg7E9RCqhGR6LUACbE
uOBvPjuuD1VLH8pBktApAybhPRqhcy1/3XOL+ueOia9tQ7dqNYzpco9UFDmACMbg
CgPgApY+rpV1IOWTe4NHEVsVa++Ax6EHzltV4TpQe2ZCbQOvg8HTSNWKy8sB0uB1
OykTTlwNiG/u/4tWcI1CUJE8kZJ6QN265WxZVYwsT5Auni1udPu+lKo+hgbMOVvo
MUykR/yhHGC6tJ6WV3rqdLFoMTXngalZegnJuOGl095nSJUgYVDtgqNe10Ym3zrX
/38wo8HMpNYWFpwp1iicdMAtA8MkJeQf/4rx9SMyT6+/MXrCe31aj2NztcIskMaL
o+Sknl+EGG8WrFw3QHLKQb1NhfPA/AtYwOIKU1FXMioq7AZT/QonOQML+lRCfI7r
CjrjrNLW3Kh/1NkBZSFO9w8staO5qCoyEyaEKI38lKxI9d5dwqsmWegEUEBHkHj+
9MqB6aCKnlB8YX0vaaPrum4H2LzNCpQyCYGvYog1ZEpwDK/R1oyYXOsp8fBcBXBt
0fYdClfkpQjXkhxIxlo1AJYZqgVnnHPBWGPZH0PhHjD6r/lGk9DZisTWNd2Mp2HN
W+R7nZaIMACLmygv0GC71Un0FcSEvJje4epf9Fi/8IETkzZy5FHzLSbKUiGEyzMg
l2aQeqyfzilezD42F5K8/8YrLEe4CWWoQSvX3PaB/kmPh1mKB2xhbrBAXS07mlUR
0PUgsdFWPGpsVwre6UgOq+aCqwHXINWghbfzB/AcV06/IkOaubZlVxF7xoZDTBwd
ImT2MfxwxXDuSHScSwT3o2odKkMhx2eVv2lQDACnqRvdrmC+C4m8F1ICPjKTHRCT
PLlhjqhV6E0hUJMrDNbZ+v8r4G6PLvgHhGtsLsnlUdzXZvzePXO+Wi0fbeZEsVpS
3ghCmJPrt9o0bhUQyMebN/XTETR1QVARVvmahupcmSa2NQ/BPof8pPW/5sf22h+X
XQYSN9V5tPO8JjkKx2gJytH61Vqeo16ZEmt8xJ9XWK7E88AK8wGhB7qxlNQo8Yrd
TfzA0GSzHrQ9ByG8H6+NUihuP3cavGG7bsQax0lD28B/Ub6haWS6gIDm7FUzkZQ4
TavPsUHTDEk1A7rkEoeDha+PzVhHrscGip91sbD8g7WapRHI6OoW/WgMt85kNVeX
O3GVUUs/3C5nvMxkb6sNa3kwm6UAN6UEly1HNwJe/QKn9jy8NSgTb7JEFPACFVuI
XsFQqerB48v4czdE3/ziwmjz7k2IXtTGo+B0+ZaJQCjo2Rjuu4X7EU2dpz05zQJ0
C9YL6SmH+PUMvH/zWzGIVHdDzP++/SDaSziEz+60Orbhh7x8l5yqGEfFjadWV7YO
OJjFPrjAIBpwQS1W/zBenhiWVCkcYOeLiOG+yzBWucTjt7u/uIsQbjQ7YPyHX94l
BByW0KSXryvGhI6rOU1JqPgY8LAVLoz1nMhC0AQelZOocOtX9/by859D/9gbObB3
8Etnl3OmN+XdzqPaXXOF1mojENbqkgBVF+D598hvnd89p2hRQNSj0uILvLWw74Ft
TpC6pUID1nNQpEvNt46C7rqEPAEvBZypjE8lgGcnYXZQ2dFOSMUe5XAE6MO666Le
ZXYmUwvST16evNg6Ez4N+ocEDleHxv+bCjorxibBzc9eGO69P7TxDTzuClwrRqxb
1zpW8cBWY9fbmLKB6szlzX9Gd7+1kBTLmglp2NhCKYmRylfnr8RimDr0J0lyDs61
gqavMFNKNnrafPgjov/L73bmGnD6dCnjsna0yBHoRifXz1TL8YC2JJBd8+h1dink
iofUA9L9DwY4aCKYATTngHvRZ5fgD9TJhxKIj5c4XXNnAcsEDPVflrkMAP1/FoHF
3m06jB2WAqWCbp6tmI7caMg3gH3WJT2fC0zbqO/HT9RpxNs7iILUSJAe8L4ejAk2
0HPUfk2iMEduMyNWsutrRnBgWxcF5MeLcFHvVBEXhbPUPqdyMj0OgtWUG1JtYSH6
Zaj3Qpse3zDoZHqm9FnbavpUnpMRiNCoCMp2rFBB4TO6Gp6XzDE044ZYp/VbUrTt
wo6n1kNOj5Yk9frMusvHSCNgirvTKopdMY9RajuC4iiMTcVkWkl+zTUQ6rI61qE8
TFBFWFEfkTGnXfgxtNq/LE22dh3Y2OU4UWWSUoWJAk188u5NalfWJdfTX/mnU64y
1gShzdhv2ZG3NgbjeZ76yYH1jDxf+MFWn9GESC4AZyKXpooJQXw0LTQXdBMmBhLg
p/888RfbiVisOC5lNPDySBk3nrg3aWVNAo5csNiU7f03+3hk5kvT5/rDiRNsJBLi
jZLtSpghciTyGjd2Bvhu5nz5dtUOSi4+QD7IDvplQo3I2ukXo1ckSXAvENqCwkLO
08zR8lDGi8ohXPQZqNAVWtPkBAkzmKLl4RXIfbh0OLv6clihg8VZtZms0/Of0YzO
QHsUgMt8En74VfCvVkXC+jGnStBH6aFEX9CTdhgAiKQ2JV4oisciMg5NT3q0nJBk
ioWCCTGY4H8Jg22jWnFtyLdYs8CNS4/aCIUl0ugA5veghWqZZWalVd++F+rbFQA8
xkGGJlRSuviFoBHq8vqqlsEd7u4YyXWDLYE5bfdhCSIaXdR25A9PdNY8R2EeDdw1
Eflsv8qzgcbmjEK31OiIDQCznQeFzgY4LtWA8csy1w7ZLNdsy0WOmYZemRSAKLBK
jdQmR37e4V+36jsjZAU/ksYyAYH423OELGjeJh3a8M0vDpC2pjrcQE35uHSTiE1R
HgT7CaYs87oHyg/ecoP0sjcTZ4KSTvZSDmC/c3SjRZxe4FMrMk7Woayh6MFG1hxw
o+yXw1OcTnH+A/oV8ozqdAZuqlp+ANlVzjvW1oKrgn0sKfltAQ13moEqGyb7h7Ci
PEloStTVzPQj+UZxGXjt81DCl3kzjI3e5RW8raqy7wY1ksKsscDNoGEqU65A/OKy
DwIy8mcdLMyYr80iGxyJWiNtsWYh6ka+kaoXEJ9IFHmC0TxpNNWZEcjV49XPoy2u
Q3R3XHdRvvjhoqjfinWhPpPxPWF9nS8I7KrRanWxi+6mDXI8LJjXOHnm6uhDt6F+
yt/eWavCUFb/5h4VdybI6zEpP8M0jQdHvkoRKNErMK7iDDNEvbHiEo4PNKxkQiKf
9mB622mKOy84t9xrsV+3z59aXbfJusX8Ff0ZOeFhGon2ydM4ZvfLKar4cBlpNEK8
UDYxXQtK1yLkecJqUvI8nEf/uGSOZmySscpmjP37qvFq+nofyiXzaQvbMwbS5YYo
wP9L/BvrW2pk5QgRRuBKy1J6NEgAmGO47tqBvHFe51Q3ZkEUlBUGTu+E1/FTGGH/
hGjUbzjO8kQwUL+IHiAlNKeCydvC5Ko3Sc1hnjoL10PfbUfnpLtjnJ/AetsW7Mu7
+oMJ5IC2kPWgv9FBIsofX9d7wUKCYmvH7wKrjCE4dyp/B6Lrq2j78NKmgEHh46IT
H7cRLGGWSafBizjNDj57Y/mN7qYX7S3DsTMJuWbfq4Eyy2eCpVOQWLBTDNlmqzWr
iznS7XkqaiVA3LzDqXtr4RAGQJgVmM0yt1FAXtqKpeiNvj3nLWIY/ifoafpL7WrE
lnOxt/BjBKneiuC5yLm6cTMJQhG8+/IYGRN0VDu1RNw6DtDmIE8uPpo19xdAhavY
HEnY23kfW2I9UhwzvDkgqF8rSFXmHcxX2WQ3lGnrYVX+sI+7M8njAp4ks6n/zON3
RCUpAGb6xBEnInTYq1NKBxem/gMBFmuSLGifx+zX/5TrmKp2AmMXdh7da5Xcztae
mS5l4BjAeoInBakUVCjSJPf+T99RWvqwZgSykfULKPwyNw1K+yg+/6+fNQ8YONWu
4cuidM6OaPNj+v0BL+he9fBOVuLL0pZM9CTAjic9rY87k0J5ICwSVwM5b6edL+Kc
lSek//oZfQTwqdhWDhRoZ5TVOFc2TQ8KF5MdAukjxu82zlg15ySXkpSWE7QUcEm3
+rBFcon92husL+I2E1cLTaNgVerD2u8fjHvjKRYD1Sqrfq4fc8imywrayVm/5O5j
C2L+UCNvr/bVSLjOVrvRNP/ybLX13TaBTtn2A6pI6ZXVmgbFOh4IBPGnq4OsGUo/
xvrzsSPvNHl4nxVUZFQFKS4DFxF0TzmdOXLrq56WB5QgpNNycWZ5flTbcse9/Uc3
nEnZSyKvveQwnfWL0osdgwmkkFZdqar4Dq2PdCnvZwwHvHKyHRz3UgtPw0SO1JH8
AESUSdvzpEpuUzWeIZTcc/LOKwmk7FEpK7eBso6bup/TOJkYNNBwstTMZGr85YeM
bUfsU2pAj69hDohPNiTpbDfx0aWDOmOBhDHVQzvlMau6d4Os2B9kn/ivJFQnqwOB
Avw2H955T9wfvqGHbMZLxjZNZsj+M4R6CjNv9VTtYe/n9YcnXQ9a7b/Fpbw4fzsl
nCRBqpnVLCgUkvKQoyMc2PpvM4WEINkCHkSggEOvLdnsC0/9bayjfWlQT/aL7jsb
JSp75n1hJmS72rf5sEmPso3Rg+STi5YTmY7nL6LgxXlxPbRO/yx4N8wNI1Jvwxra
+CQmntDec0a+4geUTkG6iRSMJ8Nnf5L8urUFn9uC10iM3Z3Tu0xhuFqedEhl6Z4d
9Zh8yFhBACZZ3qj3zx3T/20EBX4cCt7rHgyvxuZ23VpQ6KfNp9YAYO8y71djQmdI
IQNq2yZA3F8rgJpQIhkFaiyi1nQQ75RUC3ZAD3Xm+EKgmMtYlRSqY0wKkl55MHet
QBl6UjXMGBfT54GZJv1li9GcyapjjuCCGlPPSt5/q1MEnOBN54/E+ow4FULrNUMe
neQaFXz6oazFPUVJd+IfnMNiysvq9d64YkfgKOJmMdrxP0lAZODnE+nc3pe1kyOA
CqVKCmksLyYC2AVwrSZNF2HbCcB+RayDdHhQg5LPlMXf620Kjh96sR7GXPJlVJSj
HHvDLcV8P8SsdovcNTzWZk7Iy+1B2N6BhOaTV8VKmWIPCFVKpviKBW7MPqs07yIP
cUGQwWJfulMFh6ocmKFqeo7JGmdL4IpHVw3znshR6XntQm66lE49dpuZ88/fr8gI
1Xs/aR1MU9C+YjUtLHzNCFBzVOLReaByHnrTkhM+7XAUdUGsZPZnCIhaA9lIQR4t
P3Y5yCdNFDDAQjmTH9q6y5cA76SynwueSEa5IKZQY+eNWc/x+y5GUZhBA3HXIoGc
WHVo0yg2jdbqCgZC/v8G/OIDGfRWZ++TVT1aj06nH591zSokQrqowQCVQIJcl67q
ktUC7hKshougKm1TWoU8qi2xH+/4OLTJ0q96R0oMxobY4x9HCSGTUMMGmb+E81E/
tUvuHFqByS/a4enKoSSf915zwHx1bNNjyK3sfbgkZ1VRph33BC0DyukiVbsYlAnE
/RhWtytp77F6EL+tnvvadl7QEvNm3KYjLBZTrB+sWOQ/zu+AfdEgWtRXnXggnmcw
fxNL4VQMGOv07Zw/0ApLKav637DbkWVbIP8fwEDdbARK1fO/wTZmBhkrwPBHbiM+
TYt2T+CG3aQHeDPdAfoUKGMx4rS11sal0dsd1GREqsLzIIHAqnIl2uOnC05I7s2g
aq2kcMKHS5gdQlHl8F51HN5zDkbmg7fYFp64Dh9grR1TmkASpO2UtFJ+c27B5jbY
ZgVE+ZtEbHp5k78AFHcYVelLPtbzuqQ9W8xTVuhH3oUSNJOYlvWK5hVWTI6c/yqm
4GBtBZPqpqHk9cjKUK0z7zndVSQLtONBCg/8y8qKZATqf5n5pHdITTnQLUFLrX95
phgWA/ql/aevY3XVD9a3e7213QPMIBmwWtdhtlOQ2PqanBOfjHy7Fs5YzG/H2ZXP
XAdkOits9gMWPciawE0P880vLc6WKC6CY4dbYYHZkuhP1CkS8lUuoQ6iFYM1Y8z/
Vojp7EnP/T8hk0lPgg6rV6kczLTXJEUByuYT+SFiUrWjHZCFHhlyVxIfQK3R9sl8
GwZhFh++Qo6U5oKtWTRGZagCkeoYnNMxzASikDDWO2I1z2GEDvh9TOC1wdS8YlRn
dsCYDcnIm7f5GrK6FNZtty2aSO7F3Fms3oMl4dXhNskXpDNzZzUXiC/P+huXMv+6
ly5cykaFaLP6wwpoPMzKejkb2Ly4/L3tgMaKNx8Xsqcrtg7dBB2FIOWfbYLwOh04
9/ygu9NaU1nqXyyymie74h6V9I5aY1L9ze+T56jGTF4Nond/wYU+vQL10Ur+1oGS
uRBsnuwetaLjg7A8R5GulP0MVfn6EQvrz8No3U1+LASOPRqVmgbFvpu+DUKAVFiQ
hAge7+P0EYt60xiigibF9kjZk03BDJOdSQ8lwNcMNwMV+NVY961httc6eTJlIMDW
fHpTejFU42HBbBRS675Fjm8NylxUEAXe/mZ+sSokT+OQGAeSu9wT16otrh6MXNeZ
TfSdtc8zIUY1pT5PYt5ecr8jLiNCBbZm6SYPrh8Yb8am/KiZmsP/loLTCHrlrzrz
N0eANh3jUv2Sh87GK73ybKubdvQ4pV7NuA9j8hpvFhL8thH6+85VK4Qj2uBw3ref
d3MPOlHRFLqRUZi06FcN0w==
`pragma protect end_protected
