// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZH9V5jl1FJWDAAXDMD7xHi/jRDfL5vGjx8r78k8pUUEnplgZHVaPqtnkbLCq8oni
7xeq33eEHxXl74GlAs0yIyTr8NlN1PUmsIWsAAqGix1ydsl3n1IadALzbHPXLplX
/m+NhHzZ3zuTPSd+zQA4Qk6uhW7+fEPSmh/LYsBkZfQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18144)
YU4w6ScYXVBC5GG/XRvVQiNLpl6//19e1yYGYNpH4Jwy6of1x3iQ5p3yEG0YnmP0
ectwn+ooywWkMRsVeHR4jc10TtBePk/4ISLWTl2mNvIYb/24HXpHrebzYIvWODBI
cOrYtS5buUmCRQxQjei18mOu35BuKmcEme1pD3z6dZhkN+iqENrzdYFq+ZXDFuiV
nAYDPasGLOJ0jBk8Pk0Yld4RIXYTDiUYRgvarvITAFf7eAp0/1VBXo8CvV/NVWfw
qLEm8H58cSUinQC0UvOoJQa8K0hCMTSdl20aMZ5PxOPGy+uIzBUA8lQXflsIdfxS
2ferconHfah08LBQ99zGCCrPWeSqRMaTebgp4gNQsL0xwcpz6Lvnu0AJpqzISoJH
SVcxi9YfOfPb059eHtjS1z9qywn8BXuzo2wyU70qJTl6pwi8ptOecIyhQ5yo8nQn
hzzDH8Cuss2PSujqicfxZen4xXXGA18aqDwbozItcnOkOGmAUqXijfjdU7LlQzkX
kt/3r1JFrG9jOemVdpvlgYaYfZK7wHlpuenqRf7G5vGzJ1hh/NTarOev4lyej+/V
EFWC0Iu+wjfNvsoYfJjFacShN2hTNYmF2Ie53bPeLi7PQhr7OPJ5a+MFNvTE/JCt
hAic0/9w0RsgycXGaMs9s2UyJTygZH9o1d5WQ+urczvqXrG7ZT/2YCnB7DLILMea
isTBiQHcKviPs/3ey2A6Cz4aSnagCA/MCT3IXv1O3opeURF3nTgKJ6zccI8nqKCV
UHztof1mhMnklFzi4ggrRdrkdZGUGWBbpg2jle5GFzgCPpTmT/KRXDh+vbmzXojU
nqdPaDGeb/rYcZ145yoIHvuhu7HKj325sn3/SuvF1jP2A50JPr7qqu2xEHP/CFpk
w1rD9bjaAwkf8HAphUve4YNHpkaXFWgA2ZVc9jUS0wZYvMdc2bWwHT4vQp0BCi63
2agf2TotGu/lcMT9Tk3CkGBBFp4+RvviSf+QPhLVy0SQ5qc3YJ0W7XfsLZRpAbUc
KqV1dnqOMUopJRGeJNxXX0WushbeqtyQwNJR23nTRO6Gcqi30GC752/wOJiwuswV
6klr0vZ0R4z1CtQDw9EjRcoMxtzv9E6EtY98PaQUU6sDSLlE0U+3yHOGNuE40zMZ
KFznkEPQHI30PudpvZwj6LBFcJ6PciiGrtB0PiAcKySNV/qASdvap6MajSw7Q0Cl
SJaXvql6Fdhfpv8SYDY29azW9kRQubeD0MEmU3iH10mGPXYlNxFxG6+M0Lf3xlJV
QY4INgSdBDwCQJTXvHenXRsMqaIX+IfKfyEiUVjKvwOuXMHyy48eGejcAe4LJz7Q
zScjFD0RHge7u/OI7W95l4IjbwwfbEPpPY2lAgE+FcT7YBC1idU/MjhlyccgxNxe
b+8KJIfiWoBH3c78opHDTX1tv2LFIq+ELMPiMd1nooCjUFXslsvQWXP4+5BJSoTk
RAslV86FADvZaEX9Uf3IV67AKO9M/B1Opx13hLIYN3+cLrcC9pblSd0A5uBsC3fh
RxTeDG6wcKrnd//AXMrD51usWAphR3lrKDjLPtQTSa4NdzG5lINTPvyHeiDwa2pt
bijRPUuz4LxZvfErSjNXIphyj8zErboNdnqj1th4o7C1sRYldgRUCLzeTFtI2XQL
mT63YlRFLz8pwRfrzwk+cThoS278qJ/VgCuCjaMn/7Np6vEPfuoU5aAV927+SXl+
mJVP2MitSpBfKEcLq6vZDat5ODMKzktRDXfB1fJwRvBwBRtQ7SnSXyUCVFdet7S7
d7TESdudi5sYHAfqeNlIs6X6uRts3upNmwA+26Km5VK6EYfW1YUxsQd8wZLaUQvR
FaakHJGvPYeUNf4Holqw/T2s7Jd0LM/L+U30ZroUzDfQe8ipoxvKM2SC+LyLsIhC
2mjQVvnJwOpGrAxwITHaoe2KAlnOg+cjOPIA/Xj8xiSPB/EzBEW3K5Q3xl4qh7fn
0cnZkcs2XidaJHnuo2JUJV6XfuhEtuiZWz1CeWNxW0NMA6lI5RTpdy1BVne2ht5L
3ZTpVDtyMp0eb2rUYPzJNelmJnJwQ6cOtCrxjEAqoR2dMDTEC9jkXN5sP58vxo2d
CA42OhATUxcd/9oy/hhEp/EjBN/4OncxoSsD3bcr+1cKmPzIhSmFAbKPJ9/E0+7f
We06YnE2VYIkFa0pYSbzwRtOHLG0amCW2SgatkdKmjtimZ9iyUsGIyEAuf+A1UoG
1D9xZUmYTEVwo2zrM7ACFfBIXQyervtBBtveguQNga0ByNGz2E3aJP4+KZZuQIH6
0vHoyC8HzmWkWtQq1qyXFGrekyS+Qqa/gEm3qxYkbnS2Yojz1GTHzkWncu1nCYAj
CT7BbDdv1rRRQbuuQZpYSMWS+cbE+AJL1kN7RIVG+G2XaK4fVWbysZhL8Lum7TA3
KYYjsc/YiajI7k9FoOT+Q2K4f9Xv/j2sKtm256QBQ0Vh3f2huRYUI+LEGrDmy8qK
7fnCCKhNicuM59nItsyOyC0SUE//naM9Pg8a4ESzLBlkj4g8/E6tz/ps+ldkRW6/
CHyN7rcDMD5lRGKmxXEjo9pO3Wh1+MaoCIiTcqeUlfYw5HIlu0QipxpmB9ibmtve
zCFrksVHVLHOgq7FaRSqffiyMPSVHMh8zWHx4lGwYPHeYaziyTbUScnTn+BTtM3W
SSTiuq6M1oXrrCaDrnJF/1hAnltNR/QStYdAD5ZyUG74vFHOL+w4hlaFJLPzQTdK
GDp6jkjB6wYG5WkHEzb9vxeNQl4V8LShhgF6UOTtOQ86VPR5YWx4qS6feC9rpXFi
Pna2fgRqgFs7ERvT0G8kWRXSlj/+Czp52nR61EWfSju2WKzwDUuUjPu+fjFc7zwb
jaclDGbJViNr37OURotyQZyVTC+B2c/AK0dflXL6av65bGeKEnEzWMtC1T5o0vX2
6H4SlSlceDPFwHlF2pdOGmPk1m9kUXDkDtbA0PyVz7ghIKh7ixBICdhAHd7kZYtZ
vawKtyNgcecVFBG+vs9hTIo9Quwilr80S175mQt3i2LVNTJJHz8hIw1ST9o8be9C
dKlTqTxgEsGpfIoXde7I7WEpnKoA7/1TFLIKwWRjj63WDsGz8s33/bFflAwTTT14
ynSFqozMNiFuVl4FkvTyIjHgAp/zLIenhTUyw34N5WoW17OsQ5rJNTBKOnz/wyfr
yKpuOpSFW/iqz4CBxc6IzcHUOnthEeFF/6wns8g/0LdzsxDL5GLPQbJe/emPEnOz
f+jiw70kQzx+GHloYJ1BtxsZK3QqFBfS9R60vYKfAUrMhm1htrLhyZnDj9UK7ArB
VUK9EgR1vn/GsjJFISNIN4dcz9vZtQf2aifPOJcBr7fuL6cCEyO6nlpSzN2IgJFL
ylZr3jkvPHP7xD/cnn+QbVySWDfenEMVtsk8HSxWLN5wII2TG8M4Lss3V2786Nqe
tn7DHNh5SxJR8M7uq2zwMsZat7wgGWpmMu09vlKgc4oIKLVnFPIhglnOWUVSju2O
KVfAViYuOlT+AOuqtjMDugxfFu3Q4IxGmHMkAq91nRkS/vc8VUk+4TkwVBwVk7CB
6QBwNrvgj+depC/Fn9IIR3BRTJLHVWzx97RmvFscOIywpyCH3jqE3ulaiaaY4fme
Qtbtz7IWNvO7AD+/ZAjUL08qd2gN/FBEkbr56ybwxTONiVQTI99c9Q7QzImF3C9m
l4udGHR/oKzG+5GbigopCOJGKne72w8Zd/ezM8qDo3NSyfGCHExsj1K80gFQyK6R
uVhX/MbNzgO1lUPWC2m+CBlEKuWpBXhI1kgEfQuhJ5Xqks0Sar+YJZ1tltv/dguc
J6U8ESST3EvsnGgvgEtc+HulDVVJozQ9lye422rvQT6Ei+nup0oiQo6thkwWZu7h
bioyqjN632/9gYLdF93q3vn3eNCRqOoRP+saxNDHPUQNoWbIG2cGhXlY+p1b/rEX
eK8q4j/Vjy+VATXJ5jOvQapDyRPnnrG33nZLlCM6htvuvghtMs++hrZ1MGWyaLNU
soMz1xw1dH28WEBvEoIowXsT8mWl8bfSoH4emQpIFpAJ6C9wVt7B2oMTOHu3G4T+
cDisyY5w2deJPNuyuQ6r4XlOu5+TCxhT9oUbdiHEIpiStkBc+IvBviUXbDH/TjiI
1ha4sBzae8hQ4bKVlyjQd6JgDlv3Hq1pfLrzfOrWrHqjyH6HEM9upLh9ibp9sfPy
KfbxMXW66UWsdyQAL+zoJwss1a4NgdTosS7Xi3wjefFixN5gWKJEWWJbda8c3lpd
7/xiIqkSUpbcyhPF0RlrVa3+UThr1NAkM7IgmzJ2KEDUxVEMqicDojhkdcQnuKXW
4VuTSrSQZOSimMjT/yZzRgjIRWlscYrNGy+Gm+0mVUGFKIpI3AXYh/AyMYiQFo1T
QRumUALVXWeYbW53qfcQ2+tU30AUpSHTwUxg2Er2CA6eOiPGm+xKRFFGu9XS7F6o
4VPaDMiMtU8gsAqEUouBChJ/o990gLVrBRzckLBL2y/qZXsEqVPF/BcErUJYZmTG
OMXCGZfGdXNQcLp3pFEwSCLdQ0cLuAJyykq3wYdvo3Up3RKA9DqcJ5r20HkJ3ug/
QKqyfhZMT4QAm9XESjNkMHEXcORUVgnNlsutwM5xjcs9YEQDG7WPB00suIFfX3xP
/QbLv62GJgsH4xqQgUgRBXVfgInAa29flahlfnDVYB1MLww+Ke1L3ZbVMkkgz0f2
02N7o87p73PbQl4TmAYmAJiNncrGb1CzOOegbceqq7mDcJ5QyCuAQh2lr+dNOFDu
anoE1zY7H8r4J/8hHjJ+jW4jodjWWP+NHHWYHuI19qG3zvYJTE8g+BllOQqt48aO
RtFmlDicilaC3NQoB1ue+Ldifizj8vNjW1HjcCt+ZUdxcua5IKYmowANDMFThcnb
0WRWWlw/mMhIGk6FVRV+ciO7LeTH/YyBoYcVAlnF9Bqme4D+UOzmmFq17ufX6heE
7i0mYZCbMh5FeQnClWEZkA3Sz9KeBS2pi7LzoEx3/6t5OuEN2wq6p13quk0U0HOm
GBPjxTSfExTQYYXf0RAVtpisJLP28jRqJ09C6/asLoqT9bPsD70gSyEIBTTZaQ9S
Xyka2QXaIC71of7w7sMuSi2Fs3tofknpYrjkUjeXlUNykFZ2hyA6Vezsp8xUCGKT
xxu/W30323M3k9iK95HNgIY+lBOg1SOuU79A6tdTSAJO1SUNy2tADZCo69U3sQuz
as/bLY0K1E98u7RbtDK1igsKeq/NbwEDnuJ0FTUXom2K/PRuEWWm5rasde8cJMrC
7TCetfrroNU6oVpwcSu80RRWWKocED+4tASzIyvp8Br+VNGnsbwCW4feZfojtT/U
o6RSAwBx3+sUhnwB6t9ZN8f1UXnU6X+SZRIBBKi6VS+HvZ+zgw6nWL7m4KRMAuoG
6jQZ0LM+IYEU/+YdHzyBB6hXiy99yBUo4IsriFPDrRPdEAnbLCmoV7kMnYYwwGy4
/VKlZkLUrUtucmMlINjT+nVOXGOu0MP1AKRlpwY9IbZSh6924TnHXYh6ymENbaVA
7L+OM3LlN+sVKG0pcwdFY34CqQ7IBqsNZLajFzGV/CEtTTTAXwhztoHY0tjRZWsQ
6xZX5Nr30u4Z/rURQBKdoGOcjQVB5EseIWzPb9jR2XJfoumUZn1FfsIwp2zVzUIT
REC2b0/Lh07/eWl2R2En0vm7LYYJuinWTr8vrqnpVFVwCUvJx29oKlqrEaj3Oy5J
skmf1AiLtlZDpOdfduEYX8qQybo9YkYK8UOje8QHWk/ho7yBrIaz8vxG2JqlKTUD
JRVSzIVmihd/6GeEtsp8qI75QFzTs6SouZI5jiTWC2+IGX4O92JxYxeeqK1+3OKk
5fYiOoaO3ecRlKRDhXz96m6VuYthFNIgUEsJ27XhTEn1bWHwqWVpSL8MyBpl1sS/
1TH3mmeqtkBC7vSi+947fMSTD00qnkPWXGDtK6O4RkCrlRCzTb3b4mbH+i64W3rz
v2S6z5zA/U9NQ4kVoDm8pnkcdo3HYFIt6Lqq32Akqhhyajw+4vs0D8e4ewj/hfBp
+jMhDBVJhds+hv7lcK90wNSovXuhswVgPha4ME6fuT6Z0yajS7I2oaHQUM/9hYWs
kR2ZaYuanxXtb34OOt8CRBMqyzQaNNDgqRQcIEaqOqjLsnYgW/k9XSRdbIFfsW5j
R/8WrI48QV8Yg2ziypMlvng5rpcEuwtZMTefLdRvjNLZ8Wk+w8k0V77LuOY9hmCX
PEfyNffKtx1ubRdIttULua4zIlKxjnZINdbn2L8VYQcvwndAc9LS+TIi7ZdfK+M1
RrqvAYbP3xKEBsCRNu4fZbsK10CAOZ5LQD611CTlIut2DhMBri6MZ29bpKfw/OTn
V5zsMPZlJhsUr5eVgybGFPONlD+fQguOSKMIvqp9YaDbHH5m0NaRcK6sql5WhpRX
3FmHx/WP/JcrnDVvYJCwIMVM1TQMAYesUdzJc4sCwUeSW6rXuu154mJjMcQapVbb
6wo9GEJVETMChQWKbDCcHYuuvu8np6b6Pp3hOi9Hd/aO04wQIIn6oJ+LXpSHgSE0
gJcQ/3jWDLTRnIxLtupW/GvAN6BYTim8AiILoQZi8P/Mpl0VS2Rf0QiOcuSSFnG5
FVB3TNlEKTGCAjBjaiZBqyVY82pj47xhc+R2LYiDuqLxT4WgOu52zWQrk67W0y/n
1pMGGJBLExqJWhX28CeEVyA9cmeYBOvxpvrKjELiW2sUBrCSn2/DMJvXhtfRbOt+
PCrna3hK+4sLvI3bl1m1mRK7isSiHyrHhXOp6d8W6weJ0vQ8QJz8VABdZBFmzgTh
r6pDJz8u/175ycUd/aBnG6rMO/Jd//y/C26BXfXRjVJ2g/1qV8XPqk+M1H39PlDn
eZksPptxYXcBy1HjRIGuouteNnSR5Ms/PrVaK3aMpAqJIrHfO8KlMTa7inocfvk7
3pVbg8+27iI3R+HCpNjOQ9ZDmxB6UkMnJbzbih7of6Im916Y2fitIUjeE7ktNK+P
TbAa7k7jfPVqDf8lDkv+6VMAG7OjjjTRPV4EYlF7y0E2gvTqic5TtvB7ElMo9GfF
v8qvH8o+8PrRv190PVGV/R6Auh/GCo0O3asi+6AGZTwbZ6Wf6rfIQ0EYixFWG8Rt
7rMpDhfNq8BsG1P1KeTaBnx9hKwqxU540ILiaoU+Co4ASPJq+WFYWicERJHysxp3
Jsj1rwNPnMZ+jIKf/0DZxNMfL26UDIOcfOLVELiS8gY51ubSdSU8LVc6+VYi9BZ6
oPU2WlTbxqA5ZBb4vKemsCe5GO3n7MfLaZOX0oKV06jdacvKYTFMvbdvpWGxWcAc
4sY9hTuu6aHiuNO6UtktIuOuU0lty8A3oQU+QIlrRR6zeatGRGXJVIicsQEUI7Ix
7AmoSd9ALJWaD7BR+bHpao/LcD6JAliyjRwxxQiw3q7IkYJC3Cwk0WtD77mvCyLc
sWz52ja2KFKAtMnT/CIoc3/vDJUDXhvdJZ1dpOZBVT8GWaaYvBmDtqBbUganQjb0
UzD05UWNk4loW10Sdh478fGu2EXwdMlirXTAeDlILLo5pHYN4KRbRyQ7Cwj3JchT
hI8ajMSLC+WUbOxkKN1deqsuYpdBvRFp6em3T9dceRKpZS9r+hC7bp3po5NM/wxU
yb3LOwZuNTVncXnRQNdJXnqEa7ffi7zHPKo1q3IJK2VETyf8/5P+VT7G3+ZwyiWB
wKcpSps8wtjc+IVtpKtxFYlBYc6jJ2x92TCEhrnUCqGd7P+HIKwgQtdg4X/4TWPM
zLANp3VuRR1EjzfCBPBsn7kTlOXCIDj9LLeyj1NpTVC3ixII8o1kmucBdm8OhzxX
jBQE4uvGCzzZTSqwz9pEgmEfYTEeFpBEFp4EChvYOhT61ocZJErG1+/YAXf39b2I
m8PgVZchFOPIX1kdr6GR3UyCXQ8p5WTiDlAF33SDMVKGnNHrg0tJJ4DR3z29wE5D
iTqOMcB7g+bOqA7gRNlWQ5uGXMb0jSOUU1i/vr0APQ56Zvm5cp2UMoaYt7xA1pfB
QKrdvuMruQd1GqY06Z2rqbHtxE9+AASxHOijT6Ik86My5lFDMAq9k6IGS5/wUZQp
A+gD+qsosSo/YZU8D59uTz34vf6Ohw07dyclILYaiJrzwT3KFqrIGwEVp/Yn2aHn
P3SA90Ds1VNnUNNOTSW3s7iXZZkHim19VpNUQXS1PQgBHEXbztCfhIf511amWBq6
O9JZaprbglhqgihwU3CKrdjDWeTWUCHjc9udecxz/ie8FjetNaHQbDqcrE5Opdyh
VVmff+MaSogho85vrvp80pR4upT01QWqSj569K+63DojqCQnEvveEu8vsS+e84di
ZVwjUO/r+cdeV9i6FRRxESsqol/C/3RsoLa4nKGMcnz94fxNWfmE16cQSqgeBu46
BwfYKglTJiZor6LK3Hxc5Yn6L+4akH1kt2+6Anx3YPNC7gDwhhXexX65mA2e+vZ7
Ln0fL1GUjMfivp4yLXwXoqjm++2qnzL6fB22YoMv5Cyi36LU6LeRihefbSyOZ95q
OWhyQsyXZkHtfB8a0FgjvxeHRD+Toz0eg3yPvjEslYBlMUzyA1sAUzKutkTkuRQ9
98QQ1Foa8xcjuAbbvALXPIPba69Gfc6z7n+CAoaDWnrxu6VMBLbQAB8xholzyDQR
zsbG7KV+tgBBJsTwKMiFC21tYngfMOp1WphahKrtjtwD0iCOJhRvyAaxgQbZPfYW
eyOCrLARuAH5fMYCfZ2lQ5YKqiUmSzA11kzCacj0KX6HQ1sbzc7UO2sfDzTrd1TP
2P1bWumTprRNwNKMC7HyMkXclvhOFfy3cbTrZ8xaR2HUUqnDdx7FeXXTteD2I8XP
FNoVqmvbexvNdPHBkUrTsvAUCz+faJt17RmkK/CG0NOLrxzBt7V070LnWZ3eSeIB
FYTs+JZsI0GwVBT2V/sRPP65o4i77anzT2MuCSgelw3ZD+ZYXsvQiQMj37QP9AUu
Aly/AvjpCI9V4wMqHnZEPfAOs1OTlO5my/tIYz+n38RMRS0l6s86UZO7mq/AeUMj
PscfcvDkKSK/cuyyjejyZWCohVzWm/iYMDsysDlzpJEmEmfmcBazxyxXZSKNvoZU
iuieeurH4BTbQ6D+Me3+q05hNCPh00SWv0Rm7a0cdlvAJ6MW7Xh1mfL+QTX2yJbf
vBKSP1ApLsCZIiKRCWLfqFa+3Z7HywYsz9kZVXmEhRxqqS8vL1HoeeWxIjhqcXXE
102AJGoa1gnvqhaE0EH4JJLIlt0dPkJzPUY9RH+6E0vSEAWFFfds4atkwpCBf2Y/
OV9uWmvJOuJ+hKe9dYcn8YfuF3CY3b17Yam+4fIKaAvfvmFfou5PKIEa4ic68lGq
BqmgW7xy7xak4QA94W1R50/XXcL1F7EHJjydp0hxZErVuSl7Al6rdsUvOJ9EVIc6
4gyVJaSDpuorTA5tKL3czHCLj84LpJK44y75oQdqtIE6KzEwmq7isHFGiAIhqz0a
wYCagouWGmnePyUPgq5syZBZOywtiS+UWRwFdb+0zhUyflvRGSow/2yZ4iGI/R5X
Jo/8BmhXqU3YO9QFyk7s/W+SAlSZKZZWnFMgtT661FZyrCNpL8X+hKc0U1tJ8BdR
Me4C16aY7Kv9sCSGVcxmbTPR6t0xRT3Ws7FkjSZS1YyH04AqRi1bswk4vTZ4CoN5
bTTLAwDWcRxcBIk4ClyzpLtYASF42VVStHwcZNPUVcnMkAu9q7DgzVgfaYfcjmSI
cGM4JkyHgPt08phHBfUBjjRvJmprgcimm7YZlJYRbkBEPJGhG3iOQu81PbAqLol0
t23d+sgYWEOxYWtJ3besc1MJOBh+kvnOynx5oBD9BsuzvwzzLKD04zfAHDyDnfPU
lAA3pWVVnKC3FBWSBUSctH8t91zxMSs8WhgJH+5FJjrZXaccyasO3FDhL5c0pByW
hZb+VKMMk6o3JECwH5DlDOdkLaf2iScD2XzP+2AP6Lix48h0sQBioV2Whmz6f7QF
QMmUfZnR5my3B2SOCkq7WhAyiRd+fDwJmOQH5lLXdljCQL0TaLvTu5KkDJ5qvCFU
cWUV388J5mY+rOq7AhXol/2RAyHbcktSvKCacHtM+u8V4CMsJ8cvXXEc1JONPu04
JTdhdk9ZxSvVGa3BS3S12YK1TUshxO5v193PuHhayGwqvdV87Yp91TpIxv6mA75S
kYvbAxQyoLzPtOejpfdCUWmVcqjUM14T6kFol9B274s8Dgf8loSr7pacfuwqHW5h
8lpPpr3UELjCTRfuF0ZyTqgIZu0+GAYrcLlNimBI65+aMcDvmPKmL0Ui5LLAC/k8
Z4VfRBGU4ZoqgunnhHd9/KtZZdiw8VEaYHaiTTDiHjhLe3hxOR0PgC1H1CT+r+ls
qaDffQOtqmgATcu5lY26emXBfh5SnXRf9tf3lBnLl+QyLC0MH8Y0PmbRfzmNkcvN
fiU2Viem/3TFsUEkWHCdcr7PNBWsJ0pA/yhfXtv4bjnX05h7fQGeFeyGJ9aT2nST
6MN5gSdG1TLbBsEVjfY/4qNVF9ujHPu0joEtuIQnj5AK4NuP0wRhtMKJnAXumFC3
7C4NdFK4gDs3GUNIQAU02BH7W6jUkpuP7BWEaH4Fhb/9urbI2dOBddM2liDWNTxk
s1qnQdSpfNVPFu0ln6rwy/xRIJ6qu+p8rOQ2uPjF221mKlAx0wGZrsBv5PCdj5g8
JH/242QI1QHCcDRsFOkI22oMsZpv8GIAYKJFqUfEl5b8KcXEvT1l5qVlvH8iqbPl
YffWL3lVZsistAAay9z19CLLvLirBk7nV+AgH0R0wRNrAGBwUzZDm5DTW8VfcLDE
lsEsEFIYKeFIN+hia10Lec43suZNsMdia2bJfGK7NOHTQp1xWU2dwvgVB9AYwcHs
KPwhCwFPAuRZ4lvUWSDPJveVKUaQloZUnwi1ioCFEVgJAQ0n0CGMJ3vUKMvj9RpG
qp+EJhmJDzBw0Gg8kMQoSP6iyLerPlG/bEugDmkWncpY0B3cubLZRRHXKEqeTvCY
ZqEJLd4IMWf5tj1ZZGXQb9fC4Bhil56uVmnRAZ5CFdPlzLQYEw32o49PT/b1avqS
G5FyvdhQTB57GchUcao6XfNtuC945KokIvL1jn5R5z41E/1Q6V1No0MQhSWdMfKD
s20h6sEB3ivZPYv/aoLxiFfGZKntzEqWi104tYqJBMc5wOXfQcS+4BC+dLe5pKx9
7Axlr3Wih1NDxrHsIukXgTmZk7wMI0ZNl9hsW7Eof41oi7pchk+HCh62DUmXWuKi
11jzZ8DsIgMSqnysDA9murbWCFde9Z8fSvA527O6n0Y1DkhM2o1gy1qIpGilGc3c
1FcLwJvBi4XG/YJQ/9cnFHxZHpFsTSvRJ711MAp95/utDWfruJwUpKDN+UQwAFam
9ESbT40B428WgudfIIvU9rrVsbZ9zKLbeGCbZkmQSSUrVtq3bkRuqkDUcyOvN7FM
xHmCrPrYCTghxyWwcIA7htBSF/8x4G460Nd6bum1Bg3gYFAP9DTYdqeObDdcwAQm
kW1GVP1aoxDVUHckDg3+fa9MiJfIgDKX+8O0vhSV1g0Nhwu8fp+sSfkKDiZr+NLE
LeK8touneuyYIVgmBVN0FVhqSPvae9rf0WEBAl4FpDfUwNUhwM7yXCgfOuXNf1Rn
Y2cI9gRTk2WKl4xHVLwoiS33KnO5NWgT4IGErRoUe3NiXNfjASA/mQ/MyUMom4rF
lKnb1dWDgfAVaOItF+kOoBmlqrlgoQ+qFMxkJCPh6xJJ0NJ4/O0iJlWEcQAr/T32
qej3uPutXlKeBqncAuhlRDRywCT+2AL/i7WZrUE8oQfOh2Y4eMGPYyDKsAqpjJf1
CM6EMjoyMF5cgKA1Rj3kgr3FZW6rEfpdVYO/RDjiQ7RS14W1ozz+9/MfbiLOurB9
Toz4ArJ4OwwbezZh4fSEBhzDkE+AQjPdNdG2OEkC6fRa86jLUS9Fpc82ejq0ztcc
F4EJPVKCMwBqYRPR6LjQXZaRQhT06H2TapLe/8eCWLA/yz0si1SDEO5P/XZc4jxs
tYW1VktsJGTXjL1Wbwz5cAE+JEGECtQVMW7rU/mwHFIbYbe0vAvcnoWkBYmRRH6w
dvK2obviWhhw2aovrd2CeJ7KDtQtfNzUdqirafijZcBgQx29bGv1lk0ilcbtfrUH
IOG0FSYizIthz1Zgu85AuA97GGOgybN2Oq2RBdHHZBg+vymn2Rc3vxLPh0hnr9Oi
hREO7qzBLxvFBwWh6qJdZIjTXyLhOB8MKKKqm+4cHyZCswVjCIy4HHyrAwYEiU2J
SFCYdnbI5PYsCrb652kvRg98HbYc26HEg1WeE1G5GpwcsRROFYFXuZDJoWZBpnNT
cVQg9JGRpYASezUnIX5F88L08ulXzhvYo8QZ6e00zdL0CEFVzkJFc5W3nECwuyQH
YIMhMYCvkKZV4umqexd1Q0tZry8MfmSk++GGj8m2Dz3NAPFJBDNyTvjzesUS73+o
KSCtLH4bTPRS479midr0hbn+K3GQ+7UZzYQjtjCiZIOEB7tRq7KGlNK5U2Zv3jck
IyXjnMdESlTCNkfgdrX5jXrRivBg0knof/cj0tG7+qPEMVzS0BFVXt4HEuGO6b2m
0hwb73YvM4F38Omi1rhjgJC/TqqR3t0MYBfXwhfai5Iv8/l4CUEjT5AQRPKVcP2/
PVun8KgSMRGwnU+KZwnwgy5LkQQHtXEYeFO/TVreSIHly1SQueUShpP4RZsU0Jw3
7FGxB/SOkafrbJLH5fNVjYbUxiW4Yu7iN0aUZF7acwLn3XgHpOkCLjkKVJyZLeBh
f0aQJ1DSK4Ggv6fZpT0QYn97ph1gOHsbD6NACUaoU5Rx3gpinhBzRRcium/GQORj
eszgPun+6IFukcskylj5s3HnU5ijfiQwUs3Zrvi3dxABoUpOhQI1MreBB3M3UjZb
F6eV9XFlb3NKRJCDn5AnGmkj3LULPmG2w94CMU9I8dqgBqv5MJcAKUj0NzqaTWv5
kzsUgHyr5bCAdMbl24pdD9A6NvLFn5wApFS/ZgYUNCzwyz9+7oxi94xY87Fm/Vxj
bh9/7BeRwgcDojZQmX7g8rs7P6qxdnQJ77KpdDGeOoSInCQwAMcrzzDcRMUcX95l
s/t3cFwPpUdkD3W/vSjqUyhIs5ZuMWScWLDO0qk6lfKjZhYvj/SXfi7n0kvxQBSy
4nnLq6DyXkzlwMlGm8i1L+THJBiYvRoNok4OOyVvt9l5BAnTUJ0brszdNvQc3ydw
4xnCobECnn+thpE1beVIzjyaUXzhmcNvW508RD02eyGCxGtNtFBMcUi/aOYINg42
bTi/gg1QtzJwbjDxK4Y2Z+czE39FB8QTtd1RGRJ7f9S2b7kyYc53wnpye1/pFZQL
ReRP4T1IPfz07nHRmaP5pisQ9LOx+w6HRFP0q0sbQSvGKQUXOIKWom5H7l6Li3Cn
lb3v/uUnaI12Y+W2AHviGLgrYT2JN+rJEEvSqS1MNG4K8CaFr0cfBDTLKArfVrne
spEl/z5arVxRwT+3AAMBh+VQ3iPilbiRWoBp9yKqdZ5xjOAW+Jj4DVCtjwRfxduO
bHgcNUKrItG57cOeojOq9EaZhFXgW5uGK8+ZnJoONXP9Jca2tXPh81c4/4Ia5JTQ
cbmKQURxKgTfza6hOS6tI0bCWUGwbmIo3DcJgz+1QWu1sFmJ5fkJTe4mw+f2TNCY
7U90lkgMONIBFZfprQ7FL9dLja5lcNUtWu+W3AMMfXa6ahSOH7QjqeB0qFHcLgyi
+lZ0+0CucjI5j6sR7zM4msJf4YZPS2foLIdkw1hvPLGacH+ZGh5tldjReQxhQBjG
q/80iQvGvdyN5gqcThDDcTMijiBftHhzNllhWmmYvzcpH0Vym2ccGDeqhUw82SHV
OoKkdUL6MXbJnALXcq8/h8/ddUoellXPeD6KHD7Ks49MEPJOmq4RE2dAvPa5qbgO
kRDxxx2yPvzCCjbLU24NQd++ouJa1+8BJ0v52sfqzvWdA444rhoO+stqMAH1Ec2j
OUHlZDY59uNp1FYkQ2vzu7GVD4faCNDkjD5eSsvKTaexTorVwNxtVpS3nGkzphE1
fP1I3RxkTbUA2LWNgozwEbFYWUOmtiUdVUI6n4wr2viWwbOiY3f65ZHFdPiFxnkO
wpW5/mH2yZQdFi5hCY+K0+pKfaJZVfbWU1YahUuscJ9eyzlddEJ4WzOXlFtF06mj
eaw1YWFlZlW7w7d3sww7SLzqGcBX9mXgK/xtjFLdP9dQpstqJy+lZw/mnsaS6osX
hgxOT9vXN6FL7enBQ76SYPL+2n5rV6ciSzrK99I/BTa6A6HRMIMoNa0NrVmKw/XV
qgbUGJiMzSJ9AUTvqJq9N8SbK1nk4fvOucxXVRA8HiOo7ncG5Y9k5CetHxEbAKCd
2DUC5xbIbqoSJh+5xEZD+RDQoYSHIEw4JSa3OOFHP5+waLAK1kDDis3NC4Xyr42/
G9fJRULu7/QDfWtWPFdcVpnAgy4lW/B4NRqiMqjHYVxN4NubD2f0pNz64v9SXgJ8
gSDvzwCGG3QIyESBxDLusTpLxy42hsCPSPmjHd+vN7/sohEJUKUo8KNDvRGYQAFn
m7uGwQX51i6jZtZaStFD0GicOKXF2w/eTO1i32WoCgv9rcA2P8sI4P6LfuJwzpeh
+WNT2wVrxvQzF2NOnEB8b8SHqCtrmql7XiSpYlwcZZ7LJCzb8qRZmI47I3Qv/wdw
kozYRb1FpLbfz6bFE9i8S2XlmglKrfRIFOFqw4yLF2di5iJfqb6y4/wX0TBn/h9Z
9/A8i5vSDvopLTCsCo+lcwzy5bJpB5PbjobxycVURHFyK9ntwZMSSZGNzTrbJZD5
RJeuY7zSPqRlSA7KfSmVrV67O+EaMkU39R/f2cJr/aBd7wRrj4spJlUz7FbirgWx
pfgR8Oa023oO3lQF5e6W+ga0Ux8Bxy6jmLK9ZqAgM/C574qQqw+lYXhEWDFyVQqI
rKPW09LdLKHN39sPfLS/ONrJb0Y4f2UytRiM2yeD/uyHZpu5tSkv8Skc33JCKeCD
zq8l3J1gOiJV80Liglmtc8ZzDtQ+/xAJ4ZO8UX6CFXJ/s6UMSPG3qi/NZwQ6USoq
IB1IfwWwoIP5eeNsM09sbplA9AsKXCTumhSX97nurZAAyFgZNtaMD8Z377O0sppB
1XHaEuQIMHz/Q0Sjxb+oxOirNBuQJuCJwd48uy1m72VZQlVmIub/g720e652Zaiv
+6VuhbzzXfnpjVAEZJf4+eE5ALVu4JfFxzjuKymtICOO3y7/ughc4UBtU3GXqXgi
scCOl3W/nV0nmy/Zlbs4m0pbzEIf2oyWpN8yU+zjQeYms1ebaDIQMTARubIYJn/f
ssdArw8AQL1anWGXCgombB9C4K6b8tk4hFvZ7eER1kPJjZELCO82vmQ4hAkeMjFD
2Xmim+HGxXE1IUF9zSDg7U3ycRPkVswNp5UDS+xsPQ0DIkMw+lweG6MGLbVtN88j
WH8vyrNkTEdYtAi6IxtJQ1inH9tG/GcHX3kMXe7nXbMrFfbLtPUOVIhZsU4XYZpR
foz1gy0eSvonhJhQm9yZLFOO8f6qGuX6LHRx64VlQbymI3PAw47j9sCLWgFjlA3d
lgyDkjHiaUQvvh+hYWrWeW4QfZS7aIeW9bf8CQSI4GEdHI56HM3VLdHlF4nm0bgk
bvZJY5sKcD1IIvjlOcKeUrI/Khn01dKMoMzpvIoYpL8DK7wZWJ1JHma+5Yqmd1gN
TwQJXb+OuWfHf3Fn0+1kssRupmdR0HoBzX6OQtQsYwMQu3Q0NlMGMlmAAOe2v+i6
5/tRhv7j8lNfPP2HXlrPUPQvr+prSn863nURSjKWdXCWaS63n8CivOuEXVappJq2
jggu3d1TUyBNxWJ5cMhQ5vw/Qpi5BXTp7K765eQJoHM7896i6jkf9rlgQNWKJJnE
gWe4EjNhT8AV11FK0pciy2MGAkU6wcCwglyYTuHJmicuWQcJOmlvN/3N2f96v/sk
ECCUmP3K7KQvUaKKeMV1qw+kcjFqmlLJY62q8u0i3oB+I1Fz4UYCXW3Lmjoipl0L
K6hSwSL5DqPP/PuCB1y7EW0iFyiJxKdLQw9l0GOSYZ6Xyb4YAR7AAqy18Qj8C1lC
5OC4UKJEp0RJK8OQgGuvjNhykokP660ucfLlVDPjwHWIe53q8bm18IrRHAXjItax
Of83w4jGB4qdiENt4KuROqpnU5s6lrd2apDkhJgGjwkj055B6aNcw3KpMQ/TGXNQ
Pyfqaz1sySvNE6cRbVkq3LUqhfG9i2xj1ZXRdR4K1zuc3DMaTp1NRYjg2tHISW+7
U1B5YOJxfB3q9V4pJyN/+mPljQYm+3mRgQZjGMx9iCPlv66p8KO10Aw+vxHaftH1
OP+1RxiVJ335VHHk3+aGjdom4dQ5HlHaox2UYYeRe0GPiWGZRYlYV+uGlTXtmtw0
m5t0O3m6pxEeWYn6obOGVTG+l4pqNbUjvqaC0ojJFrZgFwxsLldN0iViHCWHmt6v
ifl8dv7qc9aD4eYwSp5WyAMFI32CD0YdkCmMqpBSGjoNFJErhihYWyA8j1JjYdjH
b5tE+n93U0Qk6aN2HO7QxTK/3UZbzg2MlHBMAPYxEIoHgBpxZ9KDNyu7z9rdx4QB
pNH9L20/wG8S4cMd3ZPG9G8BzGVtEG//2cAp0uFdXKA4QMrdt7pmgw6eedyIHVfl
d5/9PzmxCfeK5Rp6RS03zA3ipCheNtvZhEb/lx0hDX+KwSFnzk1niUPW4NG8Ms1W
bx6rcOsC36smmMVCp7UZ/k+xUL6Kez7iaylBo1Cb0tuS9pAy7ksGnkElicqsw1L+
WEti1/r44pfcVatj7xmzQDqQC5MmLGTdUMTChssYmVP27sdIjjlbJKqtMO4/kcLU
Rc7Mx6HbCGqmcUo52eT/dWuzJlxkgRu65ApzUZHzLTmuZmZ0AMatHzksxaneVScJ
4/BHQhxvVtGAqHUNnQ6LtmU/eFBbrxqpLkuHxa3LIQnzx+g0CNZvuH2kWoR+0P1r
XcjNnulm+f7APju3/sqF/0BjdIBHFWwzxrPeFg6BsGgIvC2MMe0pNoQU/LYtkOv8
GRlbhU/1TLDpPICFG5RgxA5yKZi7N2nMM7gaRQ5dozzGA6enk6Hsw6nw7lleatz8
L1qNPe7c+jezJFBllU9PHZHiyNByorrUJaIs6wQq7656aZ+KyclOqw/vtU9IHKnD
zEdKsnskCkPuje4FKgSuJE3Vtf8Kh3LPr/CJyRaA6fqBeA6ccf7h0hjc3o8ga1rZ
ay1X8nrCCDf9Kvx+YL1Ipexz212/zbPnZ+/ta0uNArj5+AB6QcnRrqMRcYfUujMq
rnxm/AuI1HvzoTVhZGT37yS4LuaqlMczUko5e18A3ps8A++DUOhFmSLpJ00tJ7Ux
yglhpN4zjHc3A1hclclbomMKC0rDCJ2/pmbYTtNTYppXc7CiwX2wAsf8Zf/Hdrka
IV02e9mfpb2Y2hk742NFWqywpY2DNXp6FOHgdPonmQaWBcNxXf4udIloqSi1A0rQ
w8wWY6ZzNdybnoCgDN89fFY9lo492n+Z9p/YKHTkIO89DxYIBajDd6YMfTaDmbtY
70C8F1BP8LHoyC+I1UHPKMNUDHNfcu2M6XsHqNbfxhJbtMTgiaY5o9fFImy6+Ii6
YxF7Y7o4RsnX1hKp7M6Bn55S44OagrDz8CmDjdUoJPA7vi2nmkzFQmlJk2QXYJDH
CACJZvoXvPIrOlVml2tfme6e7XKkelVTAOm0r0+b7a2nRPMO702Ty8pemZywINNK
i9P5q0ceCExQk1f8TriH7BxLYHeBvYhipLxsttgadI37JpaxDSaxtHRQA27WYEa3
KftKstHPNdKPu9yAAt5X4uXxgjd6Yv9VXBhRYjUbY/OGp/nY4NHU7TFgWjoFwxEY
c0UCnbMdaSnMrwqqhTk0dlJQo9Ny94a/bfL6ErBvHSAbGtGe4CHC5F1vYX+vurwi
e8sWtM+/bbo4hi7H3Wpyx0hBvvnmlpFYAF9GwBkxrrW/2nU/keUeiIQjF+COMPZB
nwgCZFkOuHInm1mDjezC7Yzb4ki/KmJFiLuqFhjowOwXnBamt7lzU4ERQ7b+e+Ck
aXzj5/6eK32P96LkNTQA4bPjOrao2fLv+oGkIPFbsp9eo2t6XDA0PwDcAKmxlTCF
lPOC7e8qtXEAZxN4IqbJcHH11NVgrCnsUb+loGdgMV1+4yom26Ajg6mW0+CuAPt8
CmMzm+DGxurvW8AMzbfCbIFysnEuEX5sAQzNUNtwlYRI4o3dt5048TibiKgaTLwK
wS/S31zlq6DmO6qhVyaAQnw8FQ8Xfvs/6shzhOcdyHM5Shg+MlfqHDMvqFhjcK9g
g7t2pQYjJuWtqHYRAhNb2+w4XFHiqoYlS7B01dOpoYpOHcIVcA6w10RlYjCzFFa+
bJHRA4MfY2Zy8xV40biEVIzouKzrI3pikbABWhfJSxOECq10orUnBSkuA5YoTjO3
hU8yXAOSc4CmDGrINCuHZ1FrFcQHVnGvCVllDuYnvH3FWZg1kYn5Sfnt6J4REWL0
1f9BEP2yVZ8zJKwi752QFZdS4FgRPBJQdP5YPGQTbedhm0y/GKFInCcWPtd6wU3H
NyIn88eEQY69jVlAmj41N0YEJ1TUdrPU562yof55yYJQ2MmlROo9y8jXC9LXJMB2
D6F45XdiacnKrFnTqGjSSPPEUUHzCjSzdm7gS2/4AEeEM4F/XG9jhdt6ppAsrSRJ
qCCjQr35c45tIqNnGIiMMB0Gve9TlSKxCmyEfOAvRPjMtIQpJejO6lZKHyg409Km
lCv7bU9bm070fIqreAAQAOlzyMj8C0zXdpacVhDr0w9Qf/SJ3x5PhFliggG+pGBp
s+slle13pRuuN0GBzmNlswmgPeGgOg2Qor++ggPhdUz2V5fjb88C44wSzrTqoIP1
8/cQ/+xT3xRpG2iWhQMa3MKbUvNtowN/AXK+vveEi3ie9hfEUlKn+eViBl3GKsH0
GCxdAkSYEEOU36mZDra60Vodr52KDRf6s8ROnFjtMw7n+ACGbZrSyVQFDX1D+tyv
GGIJQhCaDCmiiMKspIYDOO9ZOM5VrCVxE4WN79bMbRR6AqvR+o1iq5fCnw8V/W2O
bl1m4YBzInPRdsGkDQmhFMLJX4Qs+8GANHBhZbLGVzwCjC0TVu9OI/PgarY7b+vp
LHZKKRPaWIP4C7uUzRItkRASznVm6hjLzszz6UaNhOe7kbusm55VMfDbP8QQA8JK
kOxOSpByU27dB3EQqGhhBmsjgW53b9c8eSsFQZ9SKAa/rGpGrPT9rCKzzNsXDZN7
fGc8jcx+HrUitD7bxCKTZzm61ijmxVbHtbiU/s+6AJCGLinkB3WKqT/PoOzdU5bu
LG0+nlfXImaKeVEsXyvGy03a6953HOS6ld3X5cYrIdktcI+jqJ5G5OwAW6pUppJJ
0y8MpfJx3awy8t1qTjZUe/Br/SVM8WpQ6x7PHAor9Pv2KZLWcBeG1j2T74TYzwr6
3lXftnGgDgb+pe4GMTwEnp50ceVZafQFdv6faO+EyP01zNJ+D55mAyu1S1yPhY6E
weHvyXfsHm++o6fq4ZuDmm1rYggmpFgQZRzBODC69Wq48pab4WLYbyO6xXGKgqF5
c4NFCaHcPCG1c5ySdt6spqVx1N6JJrx42QqeWKnezbayAZI8Pz+6NeHHVnFz+H7A
c0UaReEu1mz1nm/Nb3+dU/eU/rufV56i4SI38lwapKW6l8BhQD6ETe6awb7AISM0
XqjGNXfhFF9qW+ab5Mc3gUKBOxglFc8XKSO5k+Yi6+J/olCFIeuupJwrTFbStT2C
r3nBDgBUZdhvCmLkI8GDmdTnYdqAdeZgBsNoaGraPC9HUUvJWPzm/E1QmSNmuK8v
jV2rxq0ERGTVhpVXHzfNILLb4QMkFcbR0BkYUpIz1OnuLwmW2hiYjw2WcArd6un3
EhHN2J/aWMUFisbYHNFWnBRNPaKdP/vW6/qounW41QHfoDlkkNRbDPKfl4aNGogX
+WktDawCyfxl/XZxr5JeNwHIjWEe3Y6P4YYh19c6CnQdxQqvrazQ+1x58ShICVFR
eOt7HQBJIPWNCKaNxAmsF6CZrvnXEae+Ns4Zu8zbuB873TSkkuEv4V5ZtX6wT/g6
AKnjWc9NoT0Rsl/VL2BaCvwmFRV0HhKFpFh9QDV+HMeQAtmbWDJ1APoQ9lQ39q4f
+q7GurPdFW6f0hC1YR4x6iJo7jmuAXGqVChG/4IuFSJgHBiFxPJB/Ab3GbVYFcDj
CRAei6tRisHZMWXn5tmNOeD8NI3ucfDVQxy+omwL20X/EPR31FFCwsQ7Z+g/2emY
XRP9fphm2eRVUYTkLndXLqO9Z50etr/1g/1XgW2yB5rqWmd9QygoWP7AewadSfUO
aflifhvnjfVY7yXtcIKJyOBXVAwYKSIy5lilZaxbZYbDHfDd1l62ccxicEHcJH+P
CMsK6jl6ELWvApbyh7Du60vdgO6b2vD6xWxaGq4fMbskVxZFVvXik97DLII/bYpD
yGf5mKifDajXeLgkLCEwYShT83fKr810AgODcXCzczqHjSdc/ItGFGdjTNDAjILW
H+PTY25/gbnnt+xXgP/ImypXh9qE7Fmp1LlCEnJaoxY7Zmm/clreU/BTiF0wQTml
UUDRRu8Ea0vO2i2E9EtZ8201qjv8bmKlUdAsU6LHOhk4DZ41QS7UZmYnolOIR6+i
nTKIqfbjNX2esVzsrSs7q3bW2vdBe3hFF3LTwGm7xcXiILk20xapOYqe4egKRIEh
tEtwIW9iYhhWbyqBNq48RwpLbSMUXNybBnlSmT3BFQ55iOISisabsKyAOD9Rwmov
uLn3ecN0Espw1zNSp6akrDotGeY3DiaiQcWsJNzpTUvGuXQugdOrDkUpKhVAQWpZ
J2lT034bokVZYMsRFIwgmhRCrSTF2q1pK1dhLN6VllFysSBSz0LjbhIBHP/NO48N
+dxr2pA8Z34WZXgYsA9n/lsFieIYKAIHfc0IKvCBa2QZgsRHu1AVnxe8hjWky45I
09cvnlGGwsUZV0L851j+Y+lgH2vwXdOnNeIE5yFjUK6/W3MaT+8S9oDV68DHzosp
h6KEu12yTAOadlrPy7opc4oVcvpGzXGF4yelLJP6zlDtHev9w8h/1qY9SIZgRDSq
xLlRFf5XiXiqBMv/FjUZV31ptBcQ2iPDEUrSVg4Ymor9HMtRsao8BhDnCi2aAiXA
ynbLvlgqlJ22HaZ1F6gvOPyGinXtMqzKdA6NNFBX30r+aAdb6GQQPhHZtAKgKmra
qPgWC/gDf+ngEZ5CrklXx5H7XSniZ9lDoYEiFBakmXRLOQvGR/jBCtd6DymuJp8R
O2K8XAjK8O/FE0cwlwQBN75rA/xTwADEjOSLjg3ZkUkCs4kHDUh1ka4M+jgCicDC
dINNbPqXZEMUq9ne5xUn5ksfiSLG1weCZ53BR2NXNZvohgX3sAOzqE/o7bXZVET1
sGC7/iG9EuhESrfA07idQ5pZubsR2L5t+xfSN/zDcV5PSS4+g1r6dAEz04qqcnHd
YYo1dWLmPBBRCKiUCLag5+x2mioQzeiuVdGEicMkP3LJx1lB/CwdEQ2gFJwDUTTf
VAYJy8oikUBxs6J+liQTUQViIsfAt5jLCLCAy9YuKJobN2Uoaw4cGFg6j5af3qMB
gyl108Ywq/Pz+gJknDGGLUZaqLwOcfFEb+uu7var8vnAloqxXXvXbyXqTWHXEIAV
3jaDQ8tkIg9E8d0qwk7FqWPeDvKwGA00VGzJjjep6QbI8RjOQQQ1E132cvD502Cp
syOF21EkzDtytaA1BOqBJAK9MSEG5bOqNqyqZ3UGlr0v2i3ts+uw/i7ZXOflRT+O
M5jzW8h5KszGHl716zwE3onOGSXC4O4ZSlsqbEXDl/DZJb3CulbBmIBp3x1+3Tw9
QpSueZLehzSGFeyu6fSK9gyT6aRjoIbuVt1+7LKFnCJ2moxmQKVu6NXXiSJnwKV5
134/VQdWVT3l8QvXuzPozdt2zt+AXFPw0buhm4FUO7ucxEUvwds52eGjlmbBHssL
+7H+M6DPedNPw0GOKSE7u3C94jnXnWj1dLTdabddP+LCO5DwT5/begIcr0p9f5fi
I84212L8pt/SXER6Nlwg77L9kz6EpMnjQ6xlWzDzwb5zffwFZ+jimtpMMSb8o8Xk
v1rknGDlXCgi3+K3+EjQaMLmiJ/em6g1QtdOnpLw4Y/xticL9g5ozJP4rU6vER0Q
EqQbAGeYPouva9WS2E8P3s+/sAqZxNteBl65Md/lc0s8wkU3eCe/ogRCDYZCPDJG
wu/DgjOy8wyMWyOGkNJs/ed0eI6eNRJh0yh4t0MIpIHa3LD8iwBnDB2HxzLbWxf/
QI0AFwOrVDKgipfsThbpocEo8RCl9ZnBdW8ZQlXTDLH9P1u383I4/mr7UOkN5sHA
ydg7Pqji+cs1JhMFGEPVM2M6jQeOHk7j3bvrakaPqIh8D+0/YZi0VsglzkLy1/ne
bWpElMAOD5H9JCYkdpHVH0jWpwdLqhVJWv9Sgg+gXESjyonWKqAKArZ4qjIri7gS
3Byhvw++lfJflXbHNXy7AcBwMds5B9cymx/IBwtJMdyZgaOzmEWnfHbxe8V8v9/v
nOfGIiYoCC8HK5tEHU4DRDp4+GWmVOejMhaA30ibpQPjH5joRWVVZQzHzJAQbrw3
vbvUzr2pIP1vmFCUWJnUwckPfjlVJelwPJuNyAxmgPYKXas8rlofIuT0+wOUCiHL
VOHNAwBsDqVlKglF59YgeD4akr27hjM0K5r4NfITBA26z2Fe6JRT9S1DkdviJA6B
bmUOE7gLIeeXp5wqBZfKvAOiRDthK+V00R9X5rR20cdorMUx2Yk54cDS/Sal3fLV
09Tj5mDyKbgfy3uvTpD8CohjpSAADA4ih6mFHz1uasviUYvdwGwdL24aw1VL5Cgv
gNKayqhVuaptAPo08LLWCP9p8xEuiU24eddSRnSLHQJNgBpCsze+njhWrnXg4Ru2
4aLHc6uKUzkdwVQ1Rg+P7C5DnJmoIjf8Au2jASbqhAmiO+VDwS/SCtWCnTBtpP+9
XhWHwBEkDyALr9er7FWZkW67SJsZGssyFplNqxOs6IRaX798GEAVzJao4aAg8Uy3
Hx+VDrgYHUvenP5qi7Et327OtIxSWL3n/SQQfRgArtI+XCbkP6mgbrRnLgssX+mP
c++9WueAGpPeuybQOahXiYZ/3QQVmlfwcpMZSFZULxp6t9AgBE8nM/QFS/K2Qh/e
KzQGFlHsUwpUstR1W2PG/vI1yI66PD/csE8EW/7LHUay/9wMqVoyKLHpj9MAiCIK
hvWj1pTvYuSqzsRfn/36hldcnG2kyKNuxVASvZzyd1Da8u/hD7uIqSKOuUB5Y/Ae
3vDpDDSgEyuDemyUgyTXGMRTsFf01hZBYVCTwJERtu1uYT95pT0aLaRQ18Dh+4J6
ruJZGJTPRsHWxEfCsEDw9+GzeiRqJxtWygerz3zM/jzegxh9PCO6SbK92Bkpajy7
VZDDM7HxMefpWdHIDpdMAqx58kvq++ol17V+bZUeSMPqcmgr2+fKcMou7RprWhuT
2Xj6SfPTlciPaLwMa6gO/v6ZOQP8IBal/afzLrQ92DHSZ60lHJCcTD0S5o4dMuqD
8NcsHrls1P1JPFJLrE7JKqvPDvFBLicpNEiHxLKudQgvbhYldZDzXs83z/14gq2I
L9OSvt74GsXrO9rev+XjA26J4DObH2jZYj39IRtyQla8WBSChm4jJRiNF8jeJHXu
Le5tupK4iWzVRD4lo5rfbXmJAUgHqtOFFMXYd+i9buszPRHbQn7SF03gqpmczgif
GUeDfEYu676ZdTSDGf6YsmpuhV80PqkNvG4SdUPU3vvybP4GSSFedWzDbtWTSehL
Kgcf/jKH20Dh3z/RxkTgIIvGZjSsLbmUX+ZkHAwC9nTuc1mcncweAts1XCEoBo1s
SPT0Jx7W2I0RnaZ1M2tNvRtxFWWFvuoAxLSC+Dn3HzED8K7KJgP8chuwMXowdHtU
PpiGCP52PIIAVTEpjJiGwdzwA0T6z8UshiP5SRZ1NhvIUegrMHvZO2S7Ofu5pQ1a
`pragma protect end_protected
