// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o3tjQYBTLcwVtMD0zTIeLBgjrFJ1JcVUR2cOci/vmXjTzLbsqqLQq9B4cKuHtxZe
/yYIgDMmJI4T9X9+gUCocL33PYuZ00pPcsjyROxBXEJJye6c3rYxUrwEa2kNKaa5
+wfy/F8Dwkf0QtraWpcVdE5NGkj+t7pt05aXOJiVoew=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27728)
zMG+E4VJjZXz3X8szTBylJD2E+vxpNuPLT8bVcBUed+JFTGG35BQE9zgLl+WMQok
P6jL+9qbcLDU2/eFU7Gk/Cpwq+6G9OnWPOLihSbKlKMMMeMsPuuYxFDjDOQKhpdp
l9hgnYc2LdSV4IHbeo5tTFx/1/r2JAbLSQI9doXQrFmfcmlQfsLMF4HKk28o76sf
unrvIkTki0/TU48u7/Zgf5btcW9WUnyJeA5m8riDgWQtzD3+S31SaHa9rPSHUJZI
Bhstr72LQgtqjJcts/kJUYJr90x4Zy7DJjDhZgVWI7Gi3kOZmu5VIgZj/jXfBeqn
E2Nq/rDo9okCBQXiZCKMJO1Dcv1H5v7XnlMmRPssB6NdNT/DAP5eo7/g2E0SS2u4
ysIO5s3+KeqUPCUCztivHp0miFbtcEFt1nmb5ZV+1IF8m/mLGJbWbdeY3pztmhyR
aajQ1dQdksukzot890Pt7c0n9wWQ7wM2xuyaauMs4A1rZTEick2gvQIeWUlqKKo9
JNM3xrf3cusLbbigLdZ9xUWgj2Eg+/qcOLt88db+YUjONR8hUty4Lr4XJTULXtOx
s4LAO31S/aWkP1aETwInCRGBrTE1fqdF9GKst+hNAadyL2JPB32u2W/eYLsE5p8Y
P+SwMRZIGw4In0nBH4b/Pav22k5Hsry5IKibw4ehhRCX2tBVNhndf7YlzzJkOttT
+t6hd67+dZ2yw+d1DmruuXk+ToFUAf9P4FohK7PXtnBDqrwZiTC6J8EZCnDMlNU2
jIUYiFm1u2NJWc3jZ9q4VBLbrTVKhEF75vRAVL6xHGFxgyn8z+3IRWodAgLD7pzd
rbWu2LfxxG41XFc1Rcn7tKqAWZ4B7zJz+jivtPIXl4ZMtv0nsGy52bcyH70CnRHu
28E4ECppTN7cKJfiUWPM0Oa6In6msFFSNf2pHKgz+KZ3x3OkjKLxjJJMyzOuzGQw
KniICeZ65lkYXx2ORQiqSxlOMqucKg+AslVhcd7EFfGNv1/6hiecBGPtD0LW9F1Z
UTwaHgLev5M1GMareOIOTw+0Iok18u30AbvajI3G2NA03NQX+hTA5hx2qoJmFsyU
la3N6dRZnsqqEp5W1ti1DHC9+ftnPnv5BvTz2lhktKZpSYrjCwjXPB+6b3X4Yad8
CI89jZZRPlQv6MU4tziF9rYnvyph0sTvBJa+fNhjk2RCsfTYCY15rGerWKuqzXRv
//afMVU1NPlFaPnwYXYUu7yezh7R06mrramyoOaWNE0FGPgY58qsL+DjnSpw2XYG
nxHxznJHNRHfXF5AlQSMmEr2PDexKdUQh34+9C6oLvJZnPRdkzf+vx5Oy555MonG
MfobGj5cOQHAdOwMz5f1k9uBJT170V1lIVB/PfnIPLDJWxoK5kwer05hJmxn3tgJ
TYnMZJmf8s0Z7Q5DG/Km8DyU1NWjgpfFzHu95z4AHN0xuNE7+YpFQ9jrhZYpdTD9
XMB6ao7I74GWmdJZk/CppHfrwl3VPXT3o03/7pMRDBDXb6a9RzQJlERFSnx587KV
oI6GXAUdEULbr77Yia7eoM4x2SjDGUWY3IlgiEjcmLbfH9rz3PTt4ig1MA0yFCIF
Z0sU4HPBHLKAr8GVxMP5quAAnZl4N5xyb+gvlX7sGbv86Cm+mGucvdwwonRb2k+r
78SWO7BmGrLCi+CGPRrj0Q991cZAPlh3Gx0qklnZozYzHgcDEz4KtSUYm3C3dkV4
PrNlugbgq3RmEKRsg1LOqn+y0oEamsWLEbzsCtYY+xCUrrvLD53bB+h6OFz3SULs
E44eHADxwF7J1N0eLUcS4J8i6Om5cibUYGWOlVw7L0Dy80NpwJnomczPyEI1xm8r
yTGOAnF0V2gbZTWyfMRNVKV+7j85hK1szuA8NIWO/pnYHUeo171IpLS9BNoktjqc
zYP+rq1z2iMOxcBMfheNjLVJSmVlDA42ig/L2xuGBvy/cds5tk0/vSMjWI2FA+FX
2aE6v27xecQ5VTVDoTu6MtiZ6bPEDf10JtZbF3M8ieNluPENEK1PP9+8VqmZBpxk
0adRRyEj79QRyhqnbAmtPpCZ+CQYAkBN5PTileRRx465CvKMMtudP95yxjT4lyjR
tBR0mMJFA2RWPMGDQIEe5KqaP5ENHWzROhbLIcZRg82GwDyH5w7DFsRPkH6k9f8H
uWmYbKcEz30dy6JNkEbA1MFl8wFJqm/6YpuMdukgUUjBw1HNJ4umJvhrKydVl2a+
MRRk+0TKvXKuizqdOGngQXvQWVta8zi7E3Yyx3tuWg+XaBDDFVhoL+oRXfrqdc23
5fI285dFoGccS4SQ3LTE8ZRJkgKI3vW0p+hIoszifOeh/028IsOQvwxw45EPZQCg
SLYBf4NVOWa07yte9mNdrByCGlrSPyg4rEGIJNPlz09odd0RJYbartik4EpNbSK9
89dQeoo9dkdW+SGpIgca03y5ES0a/R6YHerblEkjRfEI3QvvjRy4G1/ITfNmj6dj
oYJghwyLKdBhzxCalu43OFV+7PMcH/k9i/9VyRaaAT1rXv/RLSr2gmCCktiAx2Ih
S7mq7NMmQoyZX7J9peKGZIyFq2YFWu1HNJ9Jr0PhEOUm4gmzuFwt+WappHYCv7b8
XYwufXVpL88JFeCdHc8nfH77nSz3vK12Xb5b53FTIuwO0zBng9qJrqJRCqTjV7Ys
aopKopNCjTUaVNBDJIk+j/SutS2R0AFkcqbEX5OZNz6NmhMRFx9dmB5UTOvJtTtb
OsB/bDxAiiIEXlL8QEcYm9JOH1vJ6oi1c4JSZYAKB3nEG9wE1tvnEpTO9XDZrWkf
RL+tgsOph4BMNuNn2EnXccSryQVapROdiryxpOiazYzvWKfCbceknHBgFdhQXBy5
KRkYIpCjCjsL9zgnLhOCw5iTxf7P5yzC2lUy9ZmEJW8K/Dmd+XKMChL6abcCk5uO
i3f+ILgkK8NPd/Zp/xEGIOqAO8KC4rq6m2iCwigL/B446OJh7uCEjtzg/yjPtRW5
DH4SOw2DjRYjwIVaj+8/oTl85hQHhyA+7nZWawLeHQ/4Kf4fm3E8NJyCmlunIjRM
B1dTmvpmecFv1imSlc6DR4bUb+XRh5a+mJYGqubJ1HFGK+JCBrUaz/g8QihNqwqQ
u1RN/pMobDiqLmA+jXyrrdgGhq8Onv2i5DPvWzCCRDirYS+sTMJyZAwvLMiiAjHH
Cg/iIJfHV1sMVDtRQ94Aqk2cDC/JHt9Ez83at5eQMb9gGh01NEfJB8TWycS8bxG9
+Twz88T338cDfK620DoYRtFY0B670f7gqjo4Osjl8UA2MmYEAr52Z1D+03xjwgpr
YTsv6txTiGmYph5QEDDLJ2FcSijOk/jns8VCMmwoNk+dI0xsB5Ry5X46lOzoWESs
r4YA9SD4trmGLNhDztNO0rlW9a1xdH0E7hzWaMmX9ac9O2jWp+p+/Mr+djh3j1CG
Eu57r+h4E8T1uBI4Uf8tfNVHQfzfyyMXOapqoRYfwlUnfRJid8xT1ih+SFVVBS86
sHm60jo7fCdJWF+c/jTEgIOF9KQIg59BDeivprX31aqLTMxkHDTFoDFPGokHh5Yy
vu+L6eI+LnE73K6xvnfBBVP/Q40XaaKl94b4c08yutBraut/fJ35MmGwt6eeiT0f
DMJzFcQ1zTBo2FaYVIN0DT4j/HcLFmWaQQuqnRLiDwXFUCYbbgGI9m6v/QzkYpfk
an9tuFKIAfyUsfgUzsFz3+tUjr/6UcRROlOFyJ1nqAYrHNCZFCIvzMxbA/erv8+S
54ul7MZUenoQw43nrxHO9rYPhjQ4USeh0ortxzqoEvpfUaG0f7jmLyICUct9cozV
PyW8hR0s2LuVkN+L7j6nsYjsbD7vwMlPBZkclhYeKjcSum0q7/SpelXALb2Djzzn
GA5OBXZfAXcijbabIq9T+sVKVf+M2Rh3A1rcPM4/y2dttplTPX3Vyyisbn8ZOw6X
xIAZyI/xSvVmlJPGHC6gU9f3cFXgOSrUqKzqjJp83mzNfllcDUPPkyzEE1ucZM18
7fSSYLgZXUPjRszjaza0iOG9wEEd9I5FsdPWSVgwjXnxCt6wV1hvozemgADGpWwB
Mb2dRH4to0vYgaSHWO5GyZ9eSUihuuT74KBgkXXKW834l2fgYHm9tL93op/fpgud
uDECyPBderx8qyKQA283quQSRsNlx4eYz8ZOABX2RkiIAt4wRfSiIWyKMrnKxLFx
3RL/aMSBt9j4IlcuiSe/O9dVcfHqinpkPVbMeg3nsI0QQnJ9pWHJycH2uZ53mdbT
ye7RXrmh5QInkhvKuaFQTtwYbyYJsqa5JIZkNP2UGFfC9x3mmrVq/tJD6EO76WiD
KReM9l8WyqguVK+FKWrpunZwK1nRk4JE3/xBRvSHfjQKv3hUC4LTSs9+D+birxti
xuChKiP5HvZZ6jMzpRR8F921N9n2I9yLti+8aB8OOAvn1R8KDpnMPdeI1GdXD9eQ
0b34rimp7+rgmPd7dSCYR+XZ2ziM5TWHqjSU+fCeZlKyIz2I/4YtUJIXNwXUr/Ds
fldYBnMHPJ9O7bKcD9xw2b3aCzSbNM9rfmw10x9+K/Uv2FfM0mmzGFFmhbD7FFg8
27tJ/N0UThASmo9QXi0P2Px8pq5fnHMlV8jQLOapWrWegYRSx8BZrNMfES7EGYNV
EMlDwrcYLYhASAk0aJbLXKVDwkGOZLjnB91ZxZYews15DmlXwmXAj8AGFQTruTM0
Ju2T79xpwzkRuL9e1QfiDLM+IfJEPTz4a8D1478usf8i9kJo6uEGdZJsa0XIV/5q
SbgNqsP3yQOey6tLVDTTDu3Jmm9mSizVyjK4rhwku5H/UZZ2LifmUIuHxqXwFG1E
m1+lm+bW69LPYSnJgEGvEe1W0O2/FVQuhB9GsehSSfoiQAQxU4ggb0zhkYeQn2V/
HcdUMCnPeEoDjUdAsG222z8Vco6UuO/HY3Dn/tzgmepUsUeLTlNz7F/K3GLlQzJM
p48nqAdhJ1qAdh155CigldHz3rg/1BM0o27ry0auc3RhPOpj3NhDmpKNb04C6FjY
Xe21SQ7p6dLW2UwqjUt74oBjuS/idv0OLYIdX8FjO66Z2GLoqfOnMU9tF7jwvPTZ
sP1DZgLIX3hg4yMGbjy5sMFw9OsKFXhD95tduDTRXLJ1imMN2kwFveWQeyo7UZb6
PfHCRFB9JR8buU4c5HVjKbV66JgcgCjiYuNx2M9UdpUteJz2MaLl4EYqT3g1+QHW
u1RqobZ81w/fKvkiEiLHRHCdatdrvJNYTlVkijfzDrChPPtoK+HOnTwMhW37VcSs
Edp7wKwxfKez83hizHJVUJtpBeidfwK+SdexFM32ehHoyZrowQVOLQl2jkUtKlDK
NuDpIOtiZav7jcWdGhc3sPX5IP5qRdlqVtDaK9abTTVFy82uuHSz1xQkgxkefVnw
+XzGVyxuX6ZZSr4d8dMqx0cHwb60HQ7zk6B1jQOeYUln7mYdOvYldESNC7B9aCXK
ZvVoEOB5m0QbLwbSVFvxqjhwYNDx/odWx3a6ZsoKyEU+6xlhi2O1udMfrDOXvPCi
z0UfOeK1IV8Tt38ZWxO1OLtzIAKhcKhComOa1RSErmreKkMpFSRoFITYVr/kv91l
puK3eCv7G4YLIzHECGa9RRiE4fXqt0T6uluC8MD1MY6Mi8FBUBfKWNTfdvedUIPA
ZBxAm7/o1km73qhQES/NSpwQ2qSToJdOfVU7JXQDZItSy2+PFN1evBrQ2ENDPESK
BLInMw0wawQApB6sIaYWEoRzjQQBsaOhHdYLoPiF9DZ8J8YtmWb4I7GRjp9cM9xy
kInZTQ2Ea5W+J2rGW/oJuwto5NwoIyCvzz0jUzJBNvcCM/9u/olTh7A1khIYwdun
pzL3crNbUUthwCIDM7xHTE02DCNobs0H8zMxbBghQyxt8QFQWGJp6HdHWxOAZ1P0
6uZXfHWnqxjn7Tke1wHwAqIrt0xQBEBeB78/8HUdXA7VN4+gjOk+VIW7NasXFiBm
vXCNQipYwGq/LJyKV1U/6C1E7xtURZmFhq01yBb+8d2nhL6S1/lyTyZ0l5bBSKMv
axVHNYR7DY9E5GjEbp/fMGkjHOmQ367PkhgBrExST9CqERTtIrH++zSy8EDcxjlT
nDznbY840YwWwNG7BStX4JZJz9L/Y9LcBzr1XqiQhqIGqXb4K0bcOVENfe+IBACe
rQB/dfA/PLGje6IRTw+3MBvSyUDySHO/T9nmFRIq6O/+YHkASCCXjRx5voswx4Z5
Ecx5M7X8wT/ErfmbiZngnSHgyLPKBcvtO+sgJS18KHbttM7E/78+q7itDEIgSqc+
U/gMGPWI90wa2sJmsyhvevB/c2nepdz0wbaIrE7P0Lkit1609sZm5WRCaEzoJyK1
co8VrNZ+p2yoWkVFRFWJ53G+s714LTtETqEazEL8+gdmGYJRxLYQwF1qQNzm0IvO
akNaVyXsXw0Tpt2AohtqnWGg5Q8d9Vft0nMa6cE0mTxn4fHZoFWiy+MhWaEqWB0f
ojz+A4zMAiGmz1syzqRdpeWerdQb0rSKfjyDXiiFAEHUYsBvZsx5kv3KoWEcC54M
FUpAeS3sHKjfLFytaY4o373/hQ54L3pGEpXusCXUyZJxktF8EB5FaIcTRAwEgINj
UNiVMrFQ94w7bjLb6iQbofoVKoJ1EHKFVd5vAVQVQ6ZNsFTRAVm2bSz2pKET8OSw
z6sKuu0Sp/tTCsk1bCVIi6tSJ/uJa4XZpomzZ+hi6En6MqeOkCia/zH2Y2gAn/Zi
0OSwW8bO8YbhkMCZ7++e2EKUoE9jKkNNl6i5k8OQ5QwFNHrmMZQPcmPXsieCS75H
1iI3Zbi+AzCVdLIfgpa4UzNrwnqK2gGJ7aAvzf28QVDIfS2RW4e9p7/Wkb4kSjzR
76UIXobZ94zeNDvnLX2mElz4e4mpmDbuWXxzyuAbF8ZC+aahGnfEfomWUy1cBCx1
JjYlsanbvuo9REp5kNgP50hpxPQ3tORURSG+8jHGg46tNi4FOTwI51IySzMYmhfq
2jd941qMwMO8hQXbfJ0CZvFg9QAfPxBP3GAdMEZNEzAKrLmY/jUtBdrZZDHRrX9I
XKSSjYAq5Ucv+9ZDrwO1r4jhKMlu4ol9q7izJOzq/yIANehMn7l7U9MkDsp45aGq
2D6xiMI2HaAMiBYfZrXioZhgxSxt9pySQc/QEGDWMcR7ZPv9Ary95giqpClSzMJf
NPJa6hfLrH/etlY2F0I+6DpasgigNvyMlCc++G25G3++sP9MbDl/ZVDfCt9eqkDo
kMpdtu1YXjS1WeyaWOodz1G3znDYMj8GL4xIsB9WD4I+ctGdyG8baq9kVxnMTfYS
dQjo9198JmDvYS1epDRkJdh//XMMO0KjtZLN/pByOSjDNWtv0mQ6vzPYVsN2/x9Y
qwtILlkUMWSr0AYm2n/rp6KXdZDcJRPP9WWc5L3SXrg+VPftVn+JMWdoMOILKh6a
5eh35r0/JIudBS8Jc+672FTtH6zN/TFQaS7mrePPlVnO0GckK8ra8cMsHMBySkkY
qtdn1I0fU8rBtdr27UYI1ql9/x8RVagFRa7YFH6K4wvSNux8Vn3bR780TsHgU6bs
5snZi+J219nbVG0nOVNM3bKCRspxFzCtZesZmrhWGao4+ar+MaiEe9RS523x0MFw
i15nwKQFljud/u/XoMgVlmZLaGKqiWzKCQc6mf/nrKEjllDPK9haPRYv1uSJZMez
ST+UiGrR+dZpMwnUysMXN9QZUt5VkJ2PgMi/rD37h7a7pQsyyS6b0wWs5qFKvcVH
4PgSG5nk5R+xON1vs/aScXXyRuL4BO7XcjAE2kndHZsPMX8k5XILVJfon36TfQE4
trdJ+MiA2SEPBhYn56Jy0gSAEupZqrHgcwUq7UlWo4yAU/a7pWJMq7oLWr6OBYaq
UxpHl89Y/UUbCeRnKFGtZn4eDgQ98ZzpIJ3e5pGr+bhryHlGyKTYXjHO/X0ZAec2
oDnT6cPvSi+7g7KEAxRZToEbSeFEAp73LI/L9uf4ntymMiQNgzhEr+0R8LOrXFM6
PYOC5X7XT6CZbEeKO24VBvEAX+3UNJOIS+K6gj4Ry77lYbMvim8zqePNynCzIvSw
wE9K6CEyBXcBr9BDsk0jGnuo4r5LfJbO7zCm48tZKuJk2PI7aWVV0lxxYXs1c+Ss
xvFBERBXEXXOw7S9COi1GYiY2aylkmHMUaS815ezFvw25Bxv/zo1cLfniGv60fvV
ihYYEKdeA+phPqAr20PIlGeL1NRWuFzM6iiOdOePa48HXf7OLHx/S2cpiil3g1Sz
VfV5aS9QFmdVh8ikDMmaTGGXYXoY5Uum3B/izl1P428g2+AwsO1AF7bTfP7Q4oVm
CUGT2a2fx5VzkSCIBi0qDLfUg//js9rpW0tnquU9fJGYu/L8QQCm7F27jFbEkhD5
rWZwG5FQHEnO+eor8T3r6lXnT0LmPfK77cqyuzZRNXJqkYIGNwYh1qKI/umF3loT
n2Dp1kRsas7l9HFH2e+XKFuqPjxGrpbbd2UbmYuSBeSrDg+Y4tO/+1PV+fAGxgUO
yaz1qkT9GN5On8FNjHAZKDliH8tItXQrR8dNCfPqtIGFH7DX4WfHOrkmr1Nb+uW3
lHKbpTg0XZSEyUqO1uQpEFz5zoR8EeZsDgowv57GsEhYFVbl6HGJYSergOBWXMBl
jvzXWo/HGF7HQKAVa+5Y7a7Gtn1opZo9Ncb45WqIT8YNbnTlcG2W3ufCcXaCzXJq
nJoES/mnsyuVxo1XPLwG4eQsN0nz5Vkrc/hD5ClPdtp5sUudttxrGFWSFat/lHXm
J4/Ek6vuFRzOR576rem2lrZbnECelYP/ZwEXSufNACrUTuzCNH/MeGGJkEjoxAPa
B9zFAaggB5Iq1tn+B/PgAEfmYQPxoxYCA53X4Sl/LwaMKLDs/MZIvGmXro4UpaXD
wKQxV3NGGyWH2i0z+Ppno7SiUhnM9twYyUXCkYhZOoBNRB6BgiE3J5x10x74fmzj
m8s6zlcLgfaZqV4yCBZ5pwc48p4ucuSSr3qajGTp+ptiAsafuvrw75n1q38TDssr
ExXokY8ieFjCq/wUf3ASBhShbXAV+q8xN9lqsRZVlU6DABvHxfCCXd4B81XV2MHX
+EXkIx9brwxmLpqQViupAVSNQburLo2XHdz2XHtB1bB4IlvFHJWAEORM/Xe8u/eI
tl18R3QVFDFoMJGx3y4Cywcnjw72uxOfIDnLfwhLE7P/EbH1vjD0AtAZMPWNpqi1
Wdx5hbbZmwYSnsutnkiG4zk356V+FpiJExc6ViSKQ47KQgPwT1SHCwiYc3r0SA7w
rMgjCTnPydo0I88L6NdlKCkNXOVkjM4qGXjRNJ4uZQ1tPwigCTOO4irtXhpuWHsS
OUBpYoWKtgTCXZpTnrsoeGdvfJQmKbJoKasMzVZU5tUxbxPz4i71dQUZfAKYENKX
OJxB0rHaIa+3P7yk9nxCExlH3yNIu8FFQ/LLtnd9J4aA0wYnk2SMIlh8VVBuz9e/
36WYk9ajGPoI/+9bB1xEW8leIIA228ZScC7TC8QEhty6FGIVWHEF+CQOFAD0MliG
XTtN1cnj5EwOPasWvrR/+9HtU8dgLHCQW6QXhAxUt7WTCLZOjlOfFCKu70sS4ZkS
+ZZUZDg9cxBtDJMGyHaExIhs9f/SLfm8F+qXKV7+xl+KjL7AHvOvkOQLg81rB2yR
6+RNMv4Lvrx3IGPG40n/g8KBkg9+qFzVVFyJUgR12oNnMyhowx5GVJ/P75O63CsG
MFgSVd69OPIJi5CMTnoqxR4DH7xEi9BWfhZtB4cB8/NpVfu/IAvq6RbOHG9f7cch
Lwt2FBWwFrBgjG+R8YqdGt5oBaf8AN5YKDnGP/xFo7FOeO8cfiP/ylUI9MF0cWgt
MfLxac1XCVdWyUEU/oiOYaznr18K3y/L3NrGELqpZE7BW2edd8m8s5qh/P+QL7m6
bjhkT+uu0MNwhWV0xrNUZQV2a8Px9nyxRaND/FaPIbSb5rk8P1Rzqs2jc4MOjfdY
ZLBgWsA+x9xo5Xmn2RtSK+H38c0lpAz2z9iUDONdz4hnQmFmgmoIWwZ0xIGS8D6F
/o/cvGRvpjZq93YF52/kMNEq4eUYQOYsMmo6jWgdoVSN2vk7csV2R31IS6xj45X8
RhdKPHrM1vkEdLgN4uyxv5wSjAHEuPmDgzDnuZVMQ3m57bZ37SD+X+b8TbUJbR2/
HK/GHFzmwMmam9fHh7uovxGaYwwxcICvYID7D3OIL8SaY5DDeTHi3PWKWjrd4MsY
4/KV+TN6tjHu6aS2EJY4niXafnY2mP8vP9sVBef1JIQCVoNEsAwTV6nCVNq001Qm
rHnIoqMGEsYpiflgtV101gIUSd+q3M4t5N5FUPRORk1XkQhafadI2WXZSKO8xv9Q
RBmcHO5vbEpV2hzP5sR7uGGDATOQSl+gLcMPsJUyEnPlnroxfdiUypWdVtZeCAJm
3REWz9jsrw83nAE1ttKtXRDNpKCL0HikJ82R3edd1myUDzLWAwzQfpwpLwiixKcI
m8Kcn/+UyhvBh2yXuexfrG8XGwo/qxZ4tmDsgm5oiSVQiKpa3FmsaReOmvd8dbWE
BTW0zAAdy3FfG9TD/0yh2EfW1myjtotqgzuVFdHluTzxw10tgYcuidCQVtLL6gA9
wcBR/DZRgZTEqtGJCDJcI2F22fJTQAMz3BJXokNaGvq1JJ+HVFPlEQoag6HE79D7
AE/ahSjIV5O8j29mHWd7cZTwhIHuMro59GjbnOLF11ekeJRQ2WUfc1iNoqKXEr3C
QUzgwxQmol4wwbY3a1Vx3j9BaXKA7FBSPrutjHZPPUWjKzjf7moc2R5iCaN7uSwg
LkLzqjyf2IseIC20T7sAp5oHp2E27bFa7XfXr+xhF/r/kNy0k5wgN36gfgYxQfdK
9dVIfKEsVul+5ljegVeDSmKDh9oKGAnoWPRlwusRKGfvwM5GVmezBr42udud+9mW
QpfoFlMAuyTry4YCDcqhhGU7chlOOLFsf4mIF+xgQagQ/Yt3707Y2oNG30Wq/9Zs
v5y7sYYyYhxYqGG+yFMpfiOf+VnECkOgb6wrU0Pt+R2BSPh9R45gNLx3vTpr4cK5
Sap+z28SLlQc4QbLgWwRXgqTFoc4DHjIfZTh+ApGc9k3j8HuTHZdDgGvikHQHLic
QlDuGlTyrV1J+xVAlkZRtFFIhTj7qlZaqk0983+DAWrODJwoLHBJZb/Rci/BtPsz
4ZPHbTy87xrI0xzA7fvCUk2L8wbeZZyu0Ys/6xqbiNbx0V8uyVm40rNBoiXZMjnG
bm5AXhRxDY0YpfODpOJjC9fzfZ/QJC+QaS2+gogxt4zIQ6k6Zow2bKC4bo63q8Oy
SHmBBwPVjDsATEDTU3Dz1RTQkTLiTr2Y2EbRbjuAcAPgc/u/EiTC/97rHR7lafI+
eKesToRvVovjtgwL/jPx8mnZt9dZfTS9uN9gOD9/72buGeqVGl+EGXRlKGJj6iZe
3GrdAR6ec2kYSKZb7AldQ3Z/d9c5ZyRd9Ry1v9fUmic3NW9o4+QTfZ0Jz8UCWF+E
GHDFBLpF6cYFL+W7IVyGmylTMXfhijSDkgQidOZStUlzbS6ZZe53wo1G5J6pH9uO
LkTJXByfQ0Sfpp280+e006XwpYTCnXayxQbMUfPxDtL5o2QcR+kw0mOjaDr2TFRF
lUYgf8ed5xVA5+/sZPjypzy264EekXjPfYYsbUUapSubPWRMWoYIIPCdj1h9gQ8o
IHI+fDS6ULtsJBetdhpzO/7EWlaad1Q7TAMd8QG0U4Jjh+u6WmDwxovJqQLGmbiY
3puGuHD47GmJ5ZkUB/WqMJpV28lVJlLsyBJCnRML99vxXFjYWHEsSTXVMjILdpqf
Z6W3rTLd8HaQfNol1QaAe32bLw0ANif3jDNz+BuIlBBS/vObHd6ip8NEhc9pCf+i
FNVDUCTc/r6iHrfy/M9yP2UuUWrLhJoy7nZqs68BW6kDoI0BNrXddKTmzCCgEqI1
GXGuDYr3P9hQFEbtVueSv+MB8j0R4BCC6onr6Id5kFEs30ZTCvnE+z3fRGhV8AKs
kkdqI68JwhlYco2WuFlxcAx+CjSaW28vZCj14HJzUGljiWLPKLMRrrrYutEXpYFY
YAFEKbublVJiCZgFyN8kPNI9gfmwrBXCesvMx5NYR0zVef4EWKVcd1XzD+j2dr7Q
QIdyMyYxSCXxSfBkd3SvLEDM/CQJ1Y+gmURvhVySOByDfQ4Qo5Feje5gejFFrzgk
QaGOctBOtol0nr+GDYdIHwIEJhMP8R63LeJosm/bjL+My7mY0WNoIlCnv5WdEzVI
Os8CWcNmsZDdzRo7OTExP/kckLUL2dhVv6O+aBrZZGEpLxXd6XrlL1OX38TLi5q9
tVKpwg84jS6yk9Ch/dEsvl6cKS1m5XgciUFuw4bYOkIkXFJacAgUjm92PlycdVJA
K2HSqx8oxB0mjwkiOd//ktMkVC7CYmjcYKqZFgaM9bsfxNJgq7YaW/TIeKuQvHlA
2WI6e7wHaWfeNbxZbQxvO+JhnJvfT9ZFepJGipV3bouZwIrBo0QqD5wS7zakOU7J
dbKLk/9/gD2O5YXlHpvqcj1nICW0Zl5r1La09mRxlPGKSIxX5S5F7YwlXzG2UvlE
UvafyGCK/wc/OfzsPohT/rEKiPLsBNdsGxewq7bwrr0tDOi/eN+sPrSgEBOF1L1h
T39evqnNP2zsA/mBh2fCu6CZ6UTq3/JQs20SNSZTdW1Nv9PXFxmdZSSPN4PbSf+0
FZn8NMcLsJZqMG7sNg9GIh0l1rnwzA21DD7m572TXItkknhhtxcV9I2h1lCCVgMY
FzybBXbsE9QDhAWMTx0Jd894c+bUFSfRVeyIWWDQm5zdC+Or92aH5nij3WyqUbdl
ftmwpMCDpIcC6l8AEAiikib+mLVIm4j2PJh1YTzAEJdkNPuaF3S+ima2B3Oib9BY
Ftx65ty5eKGeulj7nxtzDu66GJcU6BNfdwSAi6omtiyOXI2JtT7+zMyCaJxfX184
mTCjjds+lTkdhNA5jTTK7f8IWyP+R+Gu8rc8jixL+7HoWC5BMxrhAz/tOGUL2yiu
ujip9Eb2dLa9gXW0aTmdKrcat6OkpHpK+yx0zKyDhBqHtFgLb+aWMtRY2OzkG4L/
YjXKy3LgBJbGPdd9P+XCxnBqenaYOLnCZoo85lnR1xG4jgNn4iq+8y0Hn8h5KKeo
lexgXm86XrGZOlgFDYEu+hv/Yu42ttPHZJ9c30Se0gRfuxC95mB4NXv83uMr8ZgA
DuyoBoEXiT/DkpLrA8nvFKYiAe34d24jcJyI3tzZoIbP2xoxTzVFMq0q2XaRHOWS
8syAuFAf6a3Y17rSs/+MNGNt/cs4CU3yt/b4DTYYEs5Hdl/O6BeJc0TkgPISeP2B
DorAV1H048yp/Xyi6qjt+nt2bHHdMH8jLnV0D5J2euY5+jy4p9F09JacEd0b3kZa
VDXQut982mh03Obn4AmRIOnrgiLt4u2bWUcqyLrw6gTUo/HKjF51NUgACuVXMTHn
TS4FIMSN9oSHVOCgnONI1rZnscVyu3E25I1gdl6bfg1Le0cxVwNZYcGyMu/38E2P
JIo0yxKJMh9nn0Cc96dTjFR6AgzxdgMYfnPPgbaXRrKUgxJDRSpyFQTdI7iUc1qA
H1SdaAwfDJGJ/q36ovvzV+YCFDngWsWgTWNNIOfGag68VHFAO9MONu0P49aRQslA
HnKusjxxHBuNTP3h8e/4IFgUOhvnf4pl3SVIz9h6crYOZa/0HMHEcS/aEkB8z19C
aJVAn9+axkWIGOeZSVEVVgrfcL+R+UlrW7vCqjZzurEZGCj3WMWWSSwT7WIlt7yx
jRvHenOAWe8lk7JR32ZEvTicX49d04su8DgqYfQfD4ibZSEomOOaDE4Xeg0Nmm0M
5GdLPxyVM68DwEFLOyuXXQaoCYIelxo1R4tMPRe8pDvtYZuDEEeqcTnEury8nQKC
Ufd2xDrW6dmoxXktkRtgCMRjDRAuiztpp0rZhYVZevSHWVs50NszZTyVpRKWDRRr
ztYyQFVz71xv89AyTF+qgtshhv+H7FbZzLev1egR6U7tN6Mtw9c9zLVXQGGRIO4F
qqa7x/9Csu/omIKL6rx8cGp1giCM+klDgaf53lU9TYSeVKMhjXQ9wRd87FpXUs9z
mwqEZCJHB4rm2TNR/Mn+9X7ntkBRs3ho8ylcYjOG6ePg5J23vUP3BptLIOGlqPRO
utxK1H1iArhmiP65LBfmMgMNdcbL7vlbcqeJgWB+Kejz5VWNIXXFhnWzWdWGElAd
106hA9U9MVswXvKFFwBlHCH5glMPlQxqvk+ToPugU4+ppYf47qtbCvRC6+eFobBZ
6M5SVDFyTSS7UOCbTrN9H8zAx6Yg7IQtedtMf282kGS6nBnQNbIqZ+BQizoNky1B
bLt+gq1abnxgXRd7H8lK/sip/ek4neaXolg7Eow3qBREGd9Q59/2m2FoFHRWdOgN
SzABsNwaSLdbYFxJh3wRhFK6BBh4XwujV4+rABUwELs7AabZP283pvlvU7/74EVA
kfaom2BQZmpGvML7+H2SAs8Y87VjfDp8+73QPx+lxSsP780M+SpPTjBSQpv3v8Dg
kf3po556xIX/PgCWFH29INnOYv63++Gn/IbCD70sWDKKL+NIjlhzaxN8HGnxRxsj
6xSQn8Zt7s5YPyHvmo9giQ9u51UPBJ9vgfy0MX6qlYEOjAkkwpSiVyy/1G8f2wxM
tD/ZL0Zq3cWQt8bzROHOl+k8QbR0R8+kO6tkG9ciy7j330Lrb8Sh6XF+2/h2Kv/Y
/vLWyr9nBq6ZRtajb1O284jM5Z9QHZGu6iwd2jNQeRjgB/e55LPBntaGL2Sdp9Vj
RGGQy1i4UlvlyJuFAJ3mNV5Pw6zAVV8EynNv7vvV0sS7fOplkW6Ozvc0ulmPONKt
GTsp1MAaWUTJEcXs6OiRDCK9oIjdaEg+F7Oo0Ze7r3cVeSrozlZNE+LYGVmyaHQb
LFNEYMCKleQI+40/VruYlvsZx+Io6a4q5jopHcEloka0glLCgI+DE/YCdy2Yt4A3
UJHH/PtzniTYZnh0gT21KxI3dcijC0bzYkYRC/9D82s5vvPFkwi7n3cBwxj0jEY6
rb1pAe39wG/ESI75CzERk1kh/nUIcwQ+xuaEIS36plO/TIq3hRhsRj/SUklyVtuf
om6YgVvvfBnHsc5GGp/2aHqdARnc0E6PbTowkGY5kC6UqLCcvON2pIIc+7kT710Q
ffHK2pPjcbswPwVzG59gZmY/ArvwE3YYDblw0EA5ZLA5CB6ZAdyBMrnTPMtxgP7Z
jgUWNxn4R2OO0rA6Nn3VDP78WRvjkKJZbubPbmmY9wTIQcGYRjQHMrmhklM5gccS
lkdzCQk3f2WkFl12GvwKgQaZPcoH1CTnVRdUwrGPKT4dTo8cTDT0ALo5L49NjqsE
Lg1PPZ3h3mCHXCJvnXVXPAz5uxfYx7iw1XFYKsqyR/v6Vf2haQQP+EwabhByfq2Q
22GmWr05iUrNUk58J1sFnhDKy6I1rd5AnKK64ux8bFfX6+XjlN2rcMZ+XqvlX2E0
vpxGdUjFvDPwP956FBzEmW/kXj/77t7plH2hJBT0HgLOi8VUnVktnhFwWmsoVtYu
Q6kIui7wBaE8/NPoMqaYUUlVY+Bqp6gBcHilG+bIwwXP11yRQHRLtzlImA+CXjG2
QH+lq6J1DBYzrbeWxhNh1E2mO+FDo0xRz7+G9olq1Ed0jWbbKHkIvBH3ta9JSW0q
urbt0aeLJ7XBEJ5yCg+yO4nyvF4ma0gTUjG2dNJpJATlLNQ53OHQfTJk+97HxWSo
FFQqCQxt1BVNjsoegoMxHOLWowHk8jZnE+YYnW4QVf31XWnJRlV5pZuLjOltIhl8
+nE+v6hi8smHuraOmvZ04jahyxPtgubD6kE6Aje1N63WISbXbAltNNmzX406CJSK
6MXLT7UAJJplMvjm3Pln7xrpP6zhaxyOii9sua1OSzex+VCoWGztvtSuhjcwv0Jt
nwMNHfyoa725uaeVxn1xc1CUVYTkciA6EmhMAzlMhddNUdxtSCsu2iusJ65yKP/j
PNYPFHUEvuLLi3DAhgheY4AcLDX+VYMubNNqYS32tU1W6GYkPTtrfLaIpIINXTlu
JuO/RHXcKViskz+fga5HqEYriAxgdC27MKbUYwgnvnENPBsvq55PuCNPhkQZlwuf
SRzFYVhjvuSmsqseRJ53OClXFUYzyzDo2/Z6tH8cGSid7qHqo+BpOAJsI8fF96t1
UR+Pg9BKSeIEUq56Eac8v0gwt8Gd/QM0e5olPgCcbMFlpsSHR572nMF0UwaZ3hwZ
22WGjIMA01HlUYR1nda34yX9ehhsqhezxQwyf10KkL2rtaJIruM4AForGbCZxh4/
4VXWTxXxFXGuBXYsQvAAM+G+BizxiJ72X+I8QPr2MgIor6okRckPlBf2mh57SBli
i3rya0SP96p3DlMOODxCrLNlkN9V4uB+dtJ4ZviaaWmGDG0lwWV87yOyPRBmjVUM
4sj+ShrjpxFWoOR1ugDXOrMZmuiNRfIOtcx5ULeeLWVVUlE9RwwjPDr1WZRT8pBf
raXpRr1dvcSsIb9oQHnbgchHndCvQEnZGoZ4QaEZ/zL/9x74mA0tiT58XPdoEIil
SXrh+GZXDaZ2BVK9y0xZr8dvRgE1L+i1Tqb4k55D9Ra51WewQAVAgmStvXGvd3y2
v9L89Cgloy5LnE6XHSkITr6qglZ8WOFg2E8yO+ukSACiIetZLFuCrZPXJmd7hVWy
dyfF+Vobg+LHaWd1OXaiN417QwP7WoEs6eIPCVxJdr1FvV4alwbziOBk8xuEIBsI
JXFQLZnG1PrDv800e3djfA0c5N4NGSS2ZQPje7+F+lDqwLWunFj8ztRlipOtJWJn
cdqPaAKoxaA5MXoT85UNIilwZUR8PpWKAlEIDrUawS+mqZEbIQqIzlv9Vx2VU1lr
dsevO115qAqWLDXm+jDQnxPslk43W7Vk1e+NRJyqYOcnEU8OaGcMTQ3ddmOUBY+o
JydHaCA0mxdg8S1RZlJovIRroXysjVKZjKkS1hHMh5IIWqQmBnWFcFlMOG/afJdt
FbWhdzVMgMLXbyzhRnXSmfmvnWvwLXzChSdt1zc3R97OFaoqiHZqbKwIWSZu28Nx
IG1MlkWcbWvVez1VgruR9SjzfKAbWZtmdD54V3ProFsSxrLGxjv1Y7dzbdBtRYtp
HMJ3E+RTUVl6httD5/vXJG8wkOQ+79jkc8r1A/YRtJh5f8qSEyp1/bWWJc2GIsul
u3fKJmMEHIpWp6tk12K/bPEh+SQHycgPj/goxkKTZD+tsUzM1n2OfukCf0z10QNG
j0aRdz4/R+d2KNy7OcYcKIn4LwuMwRyir7s34w2gauKCRf6ORQ8Ms7b6P/GNy/UJ
/ferVK/mVWhdSc9ENurUBwAJEnPsCMrMoLpR2IEefJRNi+v7nRNTWEUUHK4eX4Mh
fDUI8RAyBZQ61JGoI5wc2YS2ytK6PwG9vmVBGFcB7BYU8KPfwi6Vavz/pDoD+Q3O
ljjLp2GgwzTJDz6EmUDiQAOOk7BeWI8/5Xv9/gPcxQfdY1ciCV1lNlH6bk7yrLH6
pN9nvpia5CJ/fkIoY2iY/Ngs61bLSsp7PtNUCyQx4cS1VfaaVh5JObuFTUVjsgTa
F3o2yey3xOd+bLo575Xf+z8eWpG4a7hUnCEHer1gPAEI95q5bcCQ/00pF3No4Anu
TwNvaveQd9vNheQ/Zf1yqH8X+v3+8MRfUw9Oogyk3XSOO1hQrqKTTd1eNKFGDrdF
lZ5Ki9V4Dd+TIUw3hwWVnzsHC6cUGGdXM7r9zrLM/tqqj0icxdBNY9h3014ybcZh
eHnW2jYgJqTafLU7cZLTyfdgZ7cK9yJppX5XoMTcT6SECrUXzlrbZwX3K+ksfUs4
RUrpw0/ay+IJP6uAhPB5Jv7qfOLyAHXkhEcYTycnOyx9MYmGqYQzxJ0ZvVw/SiiT
XNIAPC6qH2/lSOsga+Gsqin4SePwUWoASuse2K3ylD+vyadTWVYrl4lUUEkjEc7V
e8LedNl8FQ3AakUpTfZn4HaYQgrk+s9Wu1R9jFtNx4ft9IeR+GpK57cxoSxRN7gO
zrGn/iKIPARFFOMqRSlW0bTjV25JlyB4CWbYlKPfkQpxKJU13xs1E98yasbu/5vj
RopwnLWxIJEK9rUFUOU2NUmw+i7KCUqQcYNhowwV3NWrot1pQshOyBs7WcLyVu0D
DXo3gx/s3zupDTk6fmFlqpyChHtoszwgaW9sq1XIHEVyRu7zzz8w7EYARd6KgLqI
jprdLnvLnHEvxP4J0D+SuKLxILlqoH2aAD++ME+6ipyK5wa4vq5CGGlZLqH3ngxv
gK8cy+QeHMluL74YECb8u5PXdxQCvtVyjkXIGaLIrOFRX8IsTQHgKV4vYAf1Eh5h
zGYgDPIAQY6jHJrf8BUPK9lhinEJOcNXukiXlAVOtlTh/hn/H+68uQSGw61i2Hvk
6hANlQhOCkmD4WY/ODa99e3B/Fy5FsCTF5ccCYk4yoIkWNKDPkqxBDuJuzaCRm04
IRjQ/xpzDwzMyNhWG3J6GZJN5ozOzbkbBVP0HFgxaVlga6U4meGeeVRHITGX+I2o
k2+2+lGuslQ/pqeFqm7RDXImpI1EZhczSZ3jqChuAGDRqM0woFtU5hkEh7tSAIYX
5BgyhUSO5OaKpIEsn0tjhmLkpJU5plmgEPeNB8SWe+EqjamC/GVGRsyiWVvo7pEX
8qzhubRECkaKKdg2NUrjLIej4++tYv/ArPXLQ+fYLF320q4Gbgjqc+r6JMaV4oL5
AvBwNz/v+VLOXd6KI19dwTmxYP/eEH2mLnSBxYx3vsXpHe7KPGb38eQXnucqQg4P
TNTnB1Pklp0cvOaNQPcPgtZJpedh1RXOJvz4/1bkh24ZgcC6Dto5VxwkP7zmjVaw
nA7AbpDH/yJZmpnzMHlxTKQRk7Sth7caFVZpOdJopqbsFRhxruZhMz5uCbtzSphw
bkvDkXMc7hGq65nKNLdGWPpWiY3RGvCatSaVAvgp3JD+unJ3EMF2vAXMTCu1Tu2a
rwFvj4RV7Qc/ig/vpTUHNwc6586lFo/1MSLvC4gZUnNvy0yYRxcIxbCxgwhdYMkE
628SOCf5K40n/K700yPfEx0xeoFMNGrfcsPqo9b5E50xjYPEDS5jQIyxMq+edVEG
6V3ANDsbCBHcRjpB5TIuwwwoUk4WGY1RWHfR1o9ZLj1xKKzEuiPT7BgfOKipIopU
N8f5JW1geXBsUyMbshSCsp01eIoi2Ie/m2KbH68AZuoIkjjsQIh4PhsM6KWNRZgO
oCtrAjdfwVnNEADnMrV9/lJAsQ7EJHQaKb6ssxYuovLEWe0BYi9tDUuM3qSMvVwL
W1h7VTrj1ZalT2P4dXmX6Eee+R/CokYDFmChnvnwrzfE2SInW4+t8eppvkYTCdZ8
6z+ChR/lQKS67u6UEbZuIbujy+USKlJHayVyzv97lH3XSvKKp28Q94fnBH+vQvmf
1CyeLr6jckiPtyRJouGQ8LpFC//4xCtMpFF/u9UBEdjRhw/bCoxSUhOfRgb17uch
nXxhbi8zK47lVJhzkELEhDM9YpugruGSyLZtRtj1q0q3KssSLikA0/gY7Y558vND
MApNO6BAa3WYJ0PmdA9Rt6PDtAmaOievidI/CUOnLUHj94fchLRmWuoFuRkFd21R
LuvijeOfQEuk77KK+tAo5NYOqA8YTLQ9/ecB/3YzFhxB7i0dun2ttDE/TbjNrewO
w4Ykde1ENknw5/nHHllpBp0FeF3sdH/iGXnNSES2pwOFRxcX4IEwmVgHmzXvaQUR
Kx1IROnfeWj1oIQFMr6YIdONlfYM5rVx29hmF28zh5HwzroddJZG2NYiJPgAzNLY
lhxejnsYwsiLjSNmg2PcMWKGrRb/jze+wkNeThx85TDGrRYi68PdXYuxhPphP/zL
5jUkfiNTJUKLe69r4VT5O8Qaz3b9FWpyYffZD00tCxHJO9IiQE2mf87CQnmymnu9
Ya4MxOOZwQqZimOKteUn7XDVy7qt7w5NSL2QDaxaXaeSRY2O/bn71WpsKNQr2HCW
F0IsksesUrdVlzhbOeEWfhla5lsWFsx1o4UL6+6tD4jXUWwaOv73XKEuAO7uuBiB
e13M4kHPIOCj/cOnXwB+mpnJALGzl1PMBQ7xXDuS7d+8EqZt3b6BsPK23iVYD3+B
gHmIMHSZqe7gRQolUnfYo3u8OzYKyhQPw3h0vlJA0KhKar0Mm0PLkTRezMvENwiB
pLeVFYJ2YWGyousuOXpYiuI1MCumRd/yYNg6WmhHbXU4NLqeSPz6srWG4bPmdms2
xvhFBqe9zYeg+6F3EcZsHy0oKY0RSbMy+F+UoT1LxnCoPBuYEe42iFf0fJi1VxcZ
n4vB0V6kYEafjXtg3r2MBmvuZj8c35mCxs2ia/ZdrlSPEqL9kF7fOD9pVZBgg6xY
r4wB4c1mfzN9Mv1udfQwyYSoia6Ybwq9S0Y5Z4U3piUYgnQoEZQ8kWrK6rkJV3JA
euRftwtmJz/k7BoDmVCTIjfnu7OV5TDSI7blkeecBCiiN4c/a3LOVhvz/nWUL9UV
dxlFqyuaZFNAyvnRSqBHEl80PmdlDbqqWWl07ClHK6p9pDMsRk/JO7sUEskgn919
gG65I6GHFAU06DNpJGkZoVinTrfVJVTAOEuD4YNmrcnI/Z6hhCOijaWKOfXf6QPa
pvljgT9UsWJC876Wq+oDb3vHaaf0N23YGA5GpRzN0Kbr6Yj1kC4KekqvLHfFY9iK
9QHxwDWDrXCuDfKp9YDseFBBAVCbpNEgkYdsGsfK680+nCTc/1jNYCQ3RfSyXV61
C1lUfrEMD2nGzl4jlOd9oV9Klhg6MhF35fmJx/Nl9Rjp5vA+mYLwdUF+yqnn/1/d
qyok/ULATmWByNL7IQZUvNu4cN7PbguYMW7j/oCFreKFxlPTwp5+JUpancmhkzlO
AmGm1Tfhw/1hxLEqjyOW8gsR6JSKn00ajpxNs9IVskLfZaO56UjTxHvBTlfYSfnY
BVVQKQ3GAkD8U6STJbHpJos7objdnL1rRoytqXL7tp1ramxvXGxhFpjPdcRhdwPW
h2SLHrPljbmOUymMZrfvqQNl3bDzjChDC1r5zvG17BTIq9eGVaeb7PyionOkbSFD
uEdpHrhQpUxBu7XlqPvVDk2tyP1ZRBnyLMtyq7QePJnmHlf+TM1tNaqBF2AnYYU4
9eJab1XF/qkE4MHbcrEcpwVcdEfAjlHv9UHzt46+EIyL72IrTFzWmLzO4Jrj+l6n
eFFFF8H2xv4Gwd/dD/pGreGte+xqOjojR6io9wTuxoMt8VOq8Qpb2KNXabXAn5Sm
oQx/ZmFTRZEaK+OUMoGVpDf1Xt7F3IvfJXhtjGsk/3+J5b3Kuc04QVB1c/KZhoBW
+tlkZSLbBgV4dOVIlNmBPIpuZvhy/BEzOGheJWRqxgm/1DMCf6onQwVOEYcmQU/A
8egI1SQrN01Wzk8v1JG26queUYb4z8IlxGaaAhYWq1FQxG1ARInqpG06phg+plfw
xsUH9YqjDrJbp493aN5Pb9AXkULqZk5mv3AofB3wD3kg5/zRr8YsvV4ax3/F4do1
BMEPXiP+hmGB/MP2mc2qJlPkcodOi8wwPFxHcIf371YAHL9ZKSVcVXYGqU06/Nr5
1Uz8Stdwf5tBOf5CwaX68Hz+1AQm1C6to7B5q+aEZBkraf5s/iOhyqqu3m8M0zbC
EzkTRyDHZ++zWlgrJu060dWmrS2ZupSMCHEI0lbIuauny/99XCB76oHhgaP2xRHz
Nv1GUvp+O4P2mca4nB6NOm5KGbYSTDbOw/xi00o3rAe1duvgwfSKTpcETnc701s1
DTt8XuCaBug96zaX6I/cD4G7WbT9zo8F77m7epymWWvKcFb03y6f0nEJgyxLWsf1
eqBR0LZzXuL5NrYxTUQTKyvlch69qhmSpidkjgwIkxEmSULcpgDIvao9MEqjcSMx
nceKrXnuHLPVrH6+mEvSx5venSHP4WNsOXuPeTFdIxXjXtUT3hEue9KCvbhrjAFb
U5f8zkNqcIFSf5gf2E7MgoT4aFs39/5n1AnYO7XVvwIRywlLVNgMu0MOF+Zv0rW5
Nc8KMw4dLxjnNZtuWpDk65vV1CuFVGSq9XYCq1Dl6+zswb6gS2KAEokPqAESU64h
wlByQwFfLl0cq2OeNIijT+oOSqPoJmq9Cw2zKw7U2CqJnBl+J9/uOb3EV+6QDXyp
enWr77veAkNT+4DoUsdwBIsKha3TO3/fkPpN+MnJew72Y1FTDjO8DinUwM0y4BhM
gJqSZjMa5T/4l3D13gKZYL3v/9B53ROGlufdr2RgXquyPMq8ZuoT5dJiUhkSwSRj
LTdfgY//1D61/vp9XmIYd9ha95zmKLzJb9CI3PVJpF8Jv3Komk8jnwWh5JmPvbed
RHC5i7P4uAGKIRJv0T8lUsE2KOdwJWygCuUTf748O3fVGZlrR17RcaEcr8T6J5I1
ZkqS+WmDxrYeUlBpx0dDx3mgIwvJIpwLvKXwhdNI8AVa4JSStWxvCbogP3hwIphp
JOm9kzqlGzZWNT2HByOLraLjGVxbQxAI95/IvvLs4sa9kQEw7UHEDPEc7J7Jud8W
J223apfl/3XzErKs53p5ODfh0MZ9d7arriIvKz/50/Pk5XiLZSbC2kdzm6C+iICN
78LMyUjlkeEumEbIlQZZF+ESAAHa5s1tPyU5Ohll4sRPoytKax+kEqPoQ8vqgYJ+
b3u4M42XpDBPe4yyC5+OIvHkGYOK3kmemeKVZA4rQ0k42iRMTwxOyY0uptzhqkTT
qdipADFER2YbInmAZdshYMQWDdBSN6vLLp/8WOENdMOazl3X6p/qvKgGlzutno7q
X6/ZkDq0qemuQHj5p+NFMI9v1/rkehfzxedLwBphnT6O7Dl1BQ/aXwllaXONQne7
WXToqTW7H7D+jc9hxJ8l8PzqdpTqe+P+/yYOG7BSvOGKnI+IiL9JaKrFJrx+WbDQ
MFb2t/J10P2H3Z2WqAQrYMMKH50DCiktYhMqo/AZKN4EXXLF3Hvl6bh5cjeTqZDH
wh3IVBUGlESI1OIglqf4l1tMABD+sZXThvhLDwP9hce8uzYePLb+Oa7iAq7Hv+pd
lKAPfb9TfsDY/NFh5YMiSEFNyiXQ5Rn0KTgB8W3RvvZ8jY98/By4MEI9nKxOQUgv
3cRF7f/nEl/Kxgw5D1awrDxDlxXbg/SlcJkJ1Q5uCrLXPswQOgezKR9VhBWmPCwi
Ckrv8ToQs3fOLClsGqelmDiMfRdRO1rauXgRC8D2uHjqJ8cnVUjkNfOPLuEnyWHP
Xiky0STg/VCBSO17SUZCgLzR/T+mG3DCXxHsr0qFmqK1HXOBKex6an7tCIt7vcLo
lWmDG+bOJUdtivJC/7jXSQtd9L+hLbUxjA0dvLJhu0BkkhCsL1s/PPkyQQSucfeW
DJEXz/DfNys00iv/XJ5OOaf8tJBBCdadFS6J52uyYm7/5qkQR10wPgmdosd09GLH
xaqCOj12wZwTiof4T6p8gn/tno/c1YEyLMNjUPWPvg0mOtNdN2kGf5jW2qS1mese
xK+wdty85GZlPbym2ZYTX16UicfHZWIR7vQ+SQBEDNtHDUVG1TqKvmZ9KMoQRGal
dgwfojAwzgT31h6jk3fYhZd1Zh7p3c1Zgr6h3nuHPGwdUHRowmL1jjy2ivBYje8C
6SaP7hZHIy/C90uXtcpneNdOFOO7Oy7iA/RaeCJBZeRQhLb1kx6XTRFzmIcPY2DG
oidYzBpvemwYbH08Iz0g1tAtgvKT/uYoxzljlhsZDlbMYweky+tdJRVwBMlHICZM
gkjgUTbdqFbJd/inBaT4SvCJfxnBy9zjRP3Q5IekwWCwCdqCeXj2ZJQlOGak5mGC
eV7fcDaEl5HvfoYLX1lv6A1WKIXUFaWd7LE8ICv5Nhxz4dnH0JB1q2l2voHkqnXV
t3cVDT6YMQIYmYaWczX6R5hCIfI63fC/Vdtu5gsOg9QxHecS1zrCayzbjB5GsoUO
FmGoBGkqpNWEKtc9bvyFnd+8TA+r45lnyENhVreDqKFrGALNHZWRDmX/eSev1W9i
LBE2fvruHx/xkmaMn5O1z/g2XHfHVAV2fhQznpBheTQKtCxwKWhFlxN9t5BwvOV1
LAvoWXWLchMX5O2OKBwvBf5arTQkQFU3mmVUKbDX/ooDRkBqVRdBDHWKkLTgg7aI
MlICako45oTuCIiuxN0sKYesFU1C5shQFDvAInRnt7f4P9Ji8q8RFWVhQtayrPa+
3Uz8T9kG+ymwBvxxyP2BC2Qtw62FjGEpJo15jivQhzF8LmaZQs2SRI9114EKjvHu
Nx4yAbg+/4C/Dk5fTPBKkxlAakz1/C0vKC7zhOc/HOlmS54/9b158QUJtr+excr0
LJJhq3dtgty+oPm62hd2gpaeuGij4ggqoijEB2Tj+wWZk9D14xfAcW9xTkfVHqpa
xMtSqvRbdMnPcHyrUOYTF5qJR13BKBRTR5oFPrBqUs0LCIUSsCaia3x2P4Q6H3zn
A3Wk8zKP7EcfSU9MWelkg+Ay7WvVDki8WEqPl4AduLAKF/qcqRmBrGOQ/SzlhFTr
BjEb9RimlvdrU6zge4v6SgoGimAu7Z/tfaZgv5iwVJPcF4oz5ANjMgP6rb16cMdL
Q6nffKUHjrvKsm17I9vSlby1GfvdC7ewueKx0yU4BM8GxH3jM5ABv0oMSm8kolFY
zsIoGvefvxpnzNId2u5hD4j9U7vcfrXTYInw7Hd3waoIi6RYNbbZ25RwO1qU/EOh
i2YVoDzjUIBhzlg448LDgNUujOH1MXhdGzV34bre2Rq+cfkpRZreO1ZLc6jzoYz2
Dg1JnlKOPgWVtauwtmCGoi4lnvMwnLRIFq5l6Cy8jOP/qn/yNvXWeLmF5mANiUcL
D348arYQAaIGsI2XBVPk79zZrPVwa8E9ZHh/GJ3IOH2DflvbmosjIOjsKrEoXYud
yHv+xNjo/ogcZ827Vfz6qEjJ9leJgpjm6zcZj4ZPVrtMOlA5KzV4JQT2OmPZ1vhN
Z4GiofNtHe+aFHKeF03Dbnyd6fGAdlgvMjQFXhPkmnQrsStXpT0nsE79MMBvGpYt
jZ065FH1XCDjKfaGAQjrPWMdyM10eUcoPU26ZBAlRzBnJ3pLq6fnvC/bpaJGGtE8
AC5CPazcfZhwbh85Ycv+vAPXxN+RXXltal2nLuChLHp0sgrC7pzqPFDgMuu1xIwr
etsl5YTBsZPcki91NLhDhFW2KVY082AHcCR8ahL+/uaqyphaLUd1/pidbzT31pXh
i1fSEcyRs1zS+mjUQ4P9Y20B6CwinILRCbU09rwaLUTfywIqW2AT20vC9nxofB3V
x03JNRomaVuq3gvwWhmurhICc7Otz7CQNJ5Xl1eXuPiLakYb2frTIzJkoG7V5VsO
bMYjSrI8ndiV8SjB6wBl4eEX34Kd9x7zPV2OZWMlmu3xlePs9CTVQGMSY+1L3/zk
evURhbtVUhVNCdkFu8GnBvFe0gZuU0CG/Odq9y6BJyTqoW/51fpk3YGm37EdSZq+
//iBjfYkaDOdo+mZzMJV1T+BL1KIpccB/ig7Y4DIAqpVsJH+xyqgokNw2xFGtCSW
jwA6TeXacJbHtxo6SS3HOkXaaOrydh63WBfcuV+xWRrNKdaOsTshCgLPOq33byza
j3OgZhHUB7FN0oc6Vm4sUNXBaZdEjXqB5JbxIjmtb/0RX5NrCfICLEqDOS8/zlPQ
umN7TkVRniX+KyVwgpIsqn5eKnO9KpH0jycZ7G0QvoaMnPpO/7lC/F/iKexcToVa
e5zLGuS/tq/kpBzFBXkFqkPKn/+XaVjf+CJTdaGoHRyZX7ty38B3k/dW2g2ZmZdj
rzX4/DPzlc2twwoLH+a7IyD8njd7hLe/trSrVJC4S+NNz0q/P/RTYFsRNZAc6ALN
nbuiFSYrU6xK8ivchIzcSi7jJtBq6oNejoTj7GBdU/wWpyL2rKEQhMELKx6kRhHE
FN6RiSfNve1ANjHjQNIVH4EL7vzJKOcpmknRG3OOY2k2twVReiLHxF7sSPEUOPSv
KYaG5pLoO5+MNHejGryGE016sS97y7qVBvLIF4SEpzV3fXbJSRe9OHrSm1nNPQKU
wqjQ4RhVLa65PuhgtzqcrCxNKTmpBHi7MQnV5XUW6S04D9FOW2ldjr2D6tw9tUMh
r+7MUSuR5aFdfXcRwaZgvs3ktnmv/1ubSichPwueYZJCZDEhqeSRkrxDg1m7J9TF
x0aIvKQyEzWEe2j4/TfSONwVonxBFulrPqzs/iJ5rvzyLrc0DcM/vzwbo+w/J/Za
9tcIDli7p9o/5UhcAQcN/yXeXhEnRZeCKN/05r+wZLZQJXePDzvFDLEb9DY6ZBmJ
aNH8KbWyq3g3AtZyZTyXV3Aj5GGs+QtbOuSyhVd2sceBkB/3N75yC6jh7E8ljYQt
zi7EjYkudKOi+UT0I0hapoEWq96BDdSUdhnLg7+fSzIImoT+Ym8YBL1/dbBXwGsv
lSpsENW6Pf04/+xztNipa3423/m7U2zS2Lh5zhXWYKZhKMn9IIG0R/l70/VIv4pw
xNsjK9D9VQHO0CtW0K+YsoFRyuzloWqtZ8hpvLM9+pFiuJzRXgxtINfiqqQFNjKB
i76vluL81nPWUD0LXv+JLhvu0FJhJ5NABox2YQOuZ2NUTu3XCztFRNjgdLQrIGMS
nz8viC13U94ihXUespprF+lQWMOWMk9RqQvfX7V7G1D4ZgYGbSREAVPSXPyoO7et
XdIiI6ITV6ntQ05hDDLMQPbChzCZYlSrFQ3TUgeGUFQkH1sXDupkliepyXsgwZ5K
VCba6pZh9yaI01fzVAfZefoiFfxkLMbSNBd7BxSWQXK48UQCyf8+CjViqDEsz4y/
k3psivpYpBegGpPACx1RQZL40O5olJnqcyy32lsII7n1tNWj0CCzivzU9zLjUA2k
RQW3ElzjtpXfKYh0IGGKEInZbAI+f7j5kf/kE6Iitnnde244iTa0WLOlkYs46ECw
MZta/zC9Glqb12X8CMas8zEljso7Ifean8QW/bocgowiEzVhwoQm8BNtp8VNo8w7
RVBqi5CpcJ2wzcYMH/WWtOrfl8YR0e2uK02LJQWPO/vimHlRJ4s7/4EnIae0xn4e
exRir9z9O1JPohl7rOypldp7x8XNYfQ5JMLWcp3KyYbIoPGEAgbw3Z3E18k43YTy
K6zvWc5t31C219KG/2eKp4+xq870kSguyURtyuWFWAf8zam4H9vaHQyXQQhy1FYR
7fyZ85ZAwUzyojh65Gy30JbzYQqMCESninGlO/CRDbbMjDQBS+EOjKNjrQetxFeG
C3GFOb39e5n9T51Ljs0jz1oUXlNeItYwuUbPChGeOhngyBU79k1ACmU+k+kJyt9C
QW/f6C/qgyAZ11rzXOkuUTSqJFylqn0Hv5L9xcdZ36pe1QVFFgcVLHzevWNR1itZ
e7sD7LodTlHto98uln4agq69KyTo9BHz7sKz3RxBiPPys2IjAgK4Lwiw3zhS7G+G
6lq57cm/tHfaR+6I/LUrTuIAnXzMYwov76cO8/DXPE67nAk9/ZOOZVY0BWkwKFM0
r/qPB8W2M44xJGTtEafu9LRt/h3GvDS9PAxwJ2M4CL1G720/ifMXzzgnBacM6Ncj
LgOeckimKkq1pokTaYpjMOxjmuc6l6YDZKgm1XCe+rnjnJB/+mZdFas2rYjDNszV
wyXNTlSYfNTp0KJui4dHYPbGfVOEFK+D/BAStcW9Pu+sjMBwIVULm0/9X/RVF8sa
uE9rZFQrHYURX9Uwu7PT5HAgtK8zkhvjch46D6HqQLAe3kyystVhkMWvHXiPCX9U
btXpJOez7m1BD4eqF6NbHJcvNS9/fXOJ0aiiSYz3mQqqmTDMMXB+tn+Jj6uUx/rZ
SRL9l1CHCr1ZP6s54YqGKpzmMC0ScVDLo+pt6MIAZsjQhm6UiYpMfwL/a3zH9+I7
mR6A50cBbSwSZ+v1dBd3cG49Brkz6UQgkryIAXJXRl+2+Cl9pYYHwn02NwwZUqaa
n6+/u1dUwe/Aq1NndTKny9aeCW5Lzv1HAB722hhZVOTiXUKIJXfxbUqBHfVSK0Hk
9z6nqr/wRBpjc6s1esm+nds6M2xQI7mQhdu8KRhIwiT0aPq6jSLvHnbPxy87ykjy
4RG6s5Lor1JijoWuB3UjHGKHZln4lGY+esmZ1NQrvKVHY6ji9H49Djn+9PFoDXQ7
RbGz81xix0PC13VNkDgN6jOxg+DBSR6qbG/yFDVLEoxVtCrYh5WLMpfJqpfPGvAo
iYMDA7Kr6g0a3wnNuBMIcrA4dzbEHt3qZKbqqjsc0A9HlxBKqbaOFORphSjEI70w
iu9StNBhbplo9LyrfTZ+VrQSJ5uOEv7dFXbvOAw+SQtF8l/AdhhY/HJWHxd895at
Cgwpg4D4aOjLbn/Vr/y225u9DRgES06rwpD+rk5sjb7ot2dPd2aRLexiCrhr+MWi
RZYkIxzhwz7bnZbuFqQYzUkLWJ1xCTR7jvhs+mBpWH7E+f4vKhQFmrRVy1IpdziE
VOmV/1nzM5aEE6vGNEYa+tpC+GxNgzKQ72TWI1PYAp73LFiRn/OrYf8sO6mLIIFv
4oRU9UnL/YWi0owms7lE5JzbtmZSaxbXOqkgcxdhSO687OhvpyNdSMl5DKco2nNy
OzZ33hofHg9kdp7zkTddHLzWJbbhiJWO4EYSavOJ4wfnQwTwe1vT/I3ci2SMeaBV
9xuF9RTzDpnwiPraxENzAAOvxJcs514kj7QVhKnNlJDVk+biAPOXtC5Pvj95yvcx
QhFSjBjUJL67AL1XP0C3IHXul+ZolFp+7MuXl6aH9Rx7YlVZtZCh2jzgBkUMUhZi
AxRisZRicGNLuhg9y/kkss9X83nRffWQaRvXHQwGavLGApoUvy0mI03tePebGZhG
vL//mm3kRG6GA8EhlAm5WIUzk7eyvFFrPWfg8YRvEf5BApyp+ea4PODXwxEGSwLt
n97wlSBxbfIGtf0x97UCne99P1AC49v8zcUB81dibpocP5CiOxm+ueSKr40mC0Fp
DOgohgu232dgHaVflbWaoy5EZLmZztHlndD5uMTKI7O4q2uiZJRozsdssaxs4avR
2A82WxlfjzrF8oTodgNA5mX2PSrysfv0fWQrmxEXEEiPC1Xq3X9/rP7yr892znPn
XVsQkt27jsVXgBGfQITVyolLIFC08L2BxQNG1flXuPtDM0SOZBZCvIBnPsSnkIah
Uu77ZC5ZYHa9IV7x5fiSPb6P0S1abz4yrMZvIqJfzRufIsz6RAMdPeJq5L3+Ks1O
nPDkLvSmNHMsmTD6z04PTNLdUIqfyNmBOj9vaJYpINSigEIrQNm+LMTIC4rwL8yZ
gmCfgI970dih3wirOvAg5qg3F8pW+bMYxDI/q+QMX0IL+A9qmBHxzejHXTEakoOl
3w4ZomYo5GfEwlefMwErc2Rmb0QIs45G1YyftbBz054GSzIl1V6aDXdo8gW3kSnd
se1E2Vmq+gZpMpL65S0u40MSN1COFsvfp4+S6QOD8E7/OPlh0J2e7zMeBFg7Miqy
+wZlEXK8Q82G5B7QryMxLyYA4UXho/EbcFPb4sZjaPYhxImZyiS6mdv+ClNqJtFb
YGC7urnOjWSKLO6aS5C24svxojKnMsvJA5ScvBbXHf8HYgNF5YJUTTtI/xpTQ3GO
L6WXXnEnoi/br59PY3gy/1kCeRYsgojilfFPZub0KNFbll/JCsvTmE+iKBzVIR2L
FHflhfonAWy8K7dZW6dHCYUXyvoB4MIAfJni5T/TljW18zcLBVsY2FV765eJJIlc
OOXEX7rzPA4YefBDQUk5tSMDjBkmC290iIkYkpAW0tizFvUoU6Xm7SLVvIEWEHl7
qt+NAyDfyGs6KcQWFmhQKmskKwYm7unzFWpUDM7k60VFccAfm71+oFMRqGYOIZvf
bvN6YdOckF1dnoZoDpbSEOf/v2Xn1mw94xGeDBVen3GVEdvFniXmL7CYGwl1dfsm
IedCBkUpZb/KYD+hMZWbjelVa2GGnv68EeTsdiJYG22qQwYAwwb1kJxSkwpn56SE
r1HFWlIW5j5jXpoaLpW/De54cHcGogsLZvcuRMxVXTiXX28o4T/UxWqR0YCzRnxy
Dx6cEddW4CRssa57cJUa60gNPV3VKJrWge1m5uL5Cu2gEfXT/EVK8p/z30R+wGU9
xaP5viG2sCmr6g0N8PmB1v31T1Yctw0pixiekW6FVQ05jyN+gl4rrgHGQImI6XRL
Dgmswvs2JsfVULM5d1t+519BDyDn8KPSKzmDB2vhDo8kZUN03g5o3pXFyYZuGxSm
YsvrXJPNDvY+WWGKH8DC5Sa/aa7wBHNsBgaaYYq7h+k09Jspa7hOwWBrV8Axtjmt
UknCOX81Jr/xS+7OogNBh/XuB4f1r+vK8mYyeL2+Bgylom83ckNHiMB1E0J5wvmz
OfE3/5tOXBc8SUmuc0rmjXl1SYvcUXQ4/H5gmeqqW8+kwHUllxBTAkHuOXtX+fKi
0mcl+HIEIgaoLYGdb5MxHBXZ46mKHWJV9cRhCurl1e4kPbWL1g4RmQR+j7AdZTwn
BCj6C9NDkoxbghne+6Ab80vaCJNVAIlsZtGGC5Y+NiLlbTO48cSSj1oPLWoHT2FM
FVMNWZYmlaKzS6hC0mfZ9MJvnZlM4AjbhO9oE/1bQMp4fPi4Q5ph5zhWnkFmIxhk
3sVCui7xCsvBbIERyIZOUFj7aouFHhfH7EGYT06DPUbz1gxYQ8emW/rVvODaFord
gvhyCc1bdoSZ7LWbcqj57ZcL1Q90OhTcdtVLuLL0cDvVDq/MSihti5it5I50OPIb
qd14jp1eoOphUiOr25SlvcS+5wpvZKeEeT7eXEWDGenV23M81DaHeLHyHZ0ewaXP
VWKTCvEkqeQhAVJqlNg//5+wyd8sWWLoCYy4uvgQCmush4A9wKOaLYbpWkH4EfZY
SuX2/FWKDwDszPBiYPf9h1eJUzjKqlXcFOMLgw64OW5BY31coPscNbLE8BZ6vuNj
U6xO4XvxA5kmElWhLE5ezsK5LdQi/ZTesa2pqPcZjjmpFlciJQGrGqPY9aalYnju
aZqRWxJJTcnfs1bOyt2WDr+gX4NADMnJiZAKEYcMpPjsXe/Z8LjE2exjYiglXYVV
KfmCwH0/BeQHx9GvG3ky8EN3STF7kCndfPQXd7CUGf9tsPU8g/dIs7oXzwuJrGoM
3BYjpBjd5jBRhigFVrQwYRgnotl28SYBnDVOw5yniCOuQErRk05RaNmbK2hU72/c
4yclEclpm5+b8dhYqBbU4/EdfmnSM7HrcRCavSWeZSr0jGuT+X96HcNWuJk2mD/Q
0KXyCRW0gKjgEMqdRpupBrJ+ePmzLpCLJimuhzl6r8Urgz9ViQBkwdUxBbKFoVkN
v9m7gwtNT5HBn1dM73sWmue2/f5lSF287dNfNNhM9bWhFwjHS8zGWRVQM5fSLqyF
0ZcEq9FXd7q/JnZDtzr7y0at1wCAhjc4hry/NbkyaOH1jOSopIZYzIGiGGqhlqUa
dmu029NvWKwiRrMFX3kTgXUlqUU1o/elkrPKyUqvr7MLkxud4roEyp7uyPndzgX8
d2v8N48bLF5fKk6OEw5KDmZavGFx1fJB7DIayEZ6wJNNOLWUMrWJtUdmK8jc/eRI
XH/UxWhdhf3alqPmdkN32wDIaDR8DPX8y+mwCkWO87GkJ/oCexK0KqJGyaQPeeHw
mqAezJuM5d1j1abuhjfDvvIln0oQpZualag19f3GLkjlAswDI5PLXC+5AK3t8yeU
Deb+Yr4RLhkvgYqHrKnCOfqlsAMHQMKmwKq9Ygox2SUf6nEFDNMpXHXFfMzgBHXj
aihFh9gQb1qDv/Bszi1cw0W1Rdk8ttLbO9/9+6+P2D8LTT4SIP8Fo8iekpILr70h
NGwoe9+f6Wtb9hHgG9dDnj+AwIEiJy4+iK/DtlrNM12rzzeOJLFwN7qYgpBT3PVL
Ge2WWOPh4gEF3slCVGRcMXVEzNNE471kYMJnxezxKwq9K2H956D1DGnisXHusKkS
oB3LXUwShAXjR+v4PuY3J/LhkdfJAEjzr4r0w5CjBfZo4MEgN13DbN/XbMbgC27c
7gMIi9pCDXYhvk1T3AcQu2/RpdPEFH+uDwDpOg66BlAHLMHnlOAVpbs5OSSWBeq9
c/bi81gdLqNFPMT0IcQO9uioli4EfnoIGedhNpKittWBcdrRJg86YuyL/4C9RUq2
HhE0tGQqR500L4+Kgm/OIwuVYbPNJ3Up6tfQUhqJ4DQxL9wh2kqj+GcxaY6ZWMjH
9VIqwuvBrTsdlObwBWWhPyNZiaETY6pYoUILjby8h1dsbTBrDB3ptMaxpol1t6hw
v/LfbvqRCXWT4mHeNrn7LCcVJzuNFpkK0hHPFl6bA5Hb/ZjTfYG70BQ8UPJs1I6t
ClKO9e8nfJY6jtfCndO9z4RPc/HdrfpW+X/w/mNSreXM12ZkMq2SLrR7gPHeFnPw
S7nXxUAn8+NT+puJGbZ563dGy0YtnoEMp/Y0YdWC/bfDY5pwCqu0mV834plWdlAt
r3l19HJFZ56y9u394xdyMrfNXc1j9M+eRoCuiLSFYybYaKz33VfKWlSo/SVZ0er7
4T8EZDNwTq35lS0MrHzn2WdFOqrxLv2RUaN/WyyzCiopUQtAhKyielNT7XtWR5zL
ZIMKKf3isWgAwzyAYk79MDpoRZhbig43K+8kBZC8i2WpESz+btZ4YbUnxwZnRGSy
6ZdqN+dxBegM4jgoAK5j5Rplz5whKRJVmL+xJjzWlIrXvBB50Cr9y7tXZ95mptxo
ohiE0VG9KKvk7L3PWQ3X8ZCpQsrK83tJi9ol9Bt5DZbo9BBSCcpXv5vQAk8USsBt
GWVB8SA7vxBiEu20H2LNlhx9Hcb67KKecokS8xM2IkGo3maKiymGCMG7aALFgRha
JNqYmnQrO7R+xwf2MwGigPSW82cuO7H2u41oI1he/AG7uPgKiq27kUFMEG8onUOp
RN7Z+kCIsDvzigjz0y0a8T+EBCpQHjjo53bhVThcMPgmd9gQN7r4TcvvjWTWy/jZ
KhF3so1PSaTNQFKE0hrmkLhxM236sgY41FHckcTTcVCbgujvje/1JmCdzplffaGU
a+gycHlU+TN7n2eQ/THdpghl0dBbMcZsAk8DFjscYFOVlXnEVovqoaWiiFR2YTvg
K6jlXzNZO22RBOvBPW5stknqu1a5K5aHpt19puJWFJ2Ysk14VE/8hd4x+2luYhHD
hNrvexr25t3UWGUeicMISUFMcAR5wFsSNi5ZL8fRpYqXtAxxx2989YTg7Rbdyr0Y
4+gQU6HA5aKo7BLTNlfIeE7SQKQCTFt3olGdx2hiLvwIaqjGZfV4hRchiriBFU1g
O+fqhQOJ4kegPGnwq1+/N1sKD93jp6VAmPDIyFNfsRfUbaGG4N+K6Qiz8x7Iq0pb
fpynXCU74SEkPr/eKORhg2i0xDloA9q+qeS2Y9IvSXar4Nb4p7YetronVoAB9Qk+
nOCKZUfcxDD2IsKwPqqly5Eh6kQgKUgC1iWB5bHsQxwqm8hJqC1GWuvU2Sbbd0yk
Ln0ZV0L0wB1UWFPTPK990Pn5GU7gy0QuNQVbT8oAYymdCqp/QwXy56bu+mHQ9+pX
Eef6ROSkw3qIDForW5LYObilIW6eP2pMw+rXsoTQy3XoRkzVqahma3tgkMnT3lVK
5DT3QsZrrwmWgb/glYNmsrNUqp3t1LqIWPVpeyU27yR+soh/K04CJM4VFu9a5T6l
JAUBI3wQbU+RhdkAgkDYZyPWxqiDUnLU0oCiHyVANQNmxJqwRi/L2TPaTSa7BcVv
y2Z3nVud5N/cYqAf1U4lcP3JdjeN3Ys8RESJnQIX+Q3TWfuCpHRdkYpPfm6WL1+C
OW/7A4+LcA/P68bdVfKto3nUDSRTXIjLnv8TE2rzn7SskK3sOcCZWtz6negI0DEy
2E9LpU3irOIlmd4BHNReqLTn4DJ5olgtkJXIm40YIq+92fJ4S9tQr/rKhAXFbIoW
/HxFOmNuOWF3fVeqG5xXJsAJ0fZ57fhLCGIBvw0xi2Dbnmd70oeAMlbjuZXvhELK
aFhkqPvhEoUhMoxrMH6aZqdGqz2frwIlJhNTuxppZZvaqxZB4xz5lQTytsGtEGVS
FNOCxMUSoMYmzwX3hBVqeLKQJKS5JinXj6n6DJNTJYxFCu6qJrQWZsG5YehDtadN
WzpJ9NwvAR/1JNpEZHcowTCKrH0by/PurJtu+6SrypVBDjYA1I08JB++d+yBk/vr
HgP8gcQYTtYEzx7xlok+4dgwecu84xNCP5DcyfugxMOQ0X31eUfD8hN8N8u85Ju9
awPIh/oPJzn0W+WQtHNqpXcMrELr84RLF1XQnemNSjHKqTPJewGvB7jTo0IUU3hL
8aY4CQTV3ismi/fZ31BdiZevXixLuFX3DooGrgP3Iw95oiLFSIDxO0R+cVeTexUy
kQKXsx1KwGXz8imLMYRp4UHhPp4PTRGXPykP0Hz1nwVQVR5zHons72+jCqjMEh5Z
j4gaJYjOQkb/VvLVR3H8K8SmUVEbeHyX51IawTyaTBSDbDLX5Asbx/3FwU8zW4Mr
vU8dDwNjHKdjrzGISohhIQSrnv13joMTVBbQ1jioKhjXig6M7LNWQNLu5+KtHS2A
qEh7B4bna5dbRMlFQfRUblDG2VRSvARJ+8wRVHvyrHOx3sleoGq3K7sHMmjgDbBA
nyokA8vA9tUTOglcQgxJ7aTcx5r5Ca+Vp11EDD0nJF8RcsnCYapySkXi8Xj5crqy
vIj62jsSFlkMA2fp7uuIot6YNM+1Sy3uj3AnZ5CyVYakBWUh3UnHsUEMlLq5dzUn
vXKJaBcE/jotCwXNgilQWpZ2CizjhJaRCPRJ+8l79M/nbtkFeQ+NT9JeAyDoCY32
S0twZZGM8Bu0LBMpmI/WP4Z4H9B12xP929glUvrHpU1kuzO/2sKYJooFbS1NB/Hs
/n30DpVHe02RfEldVVOhr8mN7FFb35oKZeusegPsCNC5+pxIeKN5zOYr8/PCKBaV
e9tg2ygtOvFKNzv0gqmNnEOeM/TU0plFe1BXH6vPIHXT9x5cHj7IU38rjOTBCvHO
vWKcfBzxNXj2uXBPTzIsu1XXf6PhPBCTTEBy6kU1ZhODJsrboRlkgk+Gkbdtn66D
RdCp7cVLr9jJwtKLOLH9hNYbSIRSx5Nk9m+BKK2pFsg0bxTqVhg+TTVfxVynxk4p
yNapexRcqU1ZKwCFGefQ5fI5/08/TB0Pf8dGyz/5k/E6axmkPD+xUt5+cu80NAAF
cghiesdEajAf04KGnkBOyvAKZdnqVdK1nYT9jPTczTzhBeF3W+cjNNkDEvNGOw1e
rDQKWmo0KHPPCoDmXKwr/OryfeY7F7qH+yNbKt/XdDegeiLsPhnBrY7lrsHkikUe
n871GdGuzmcjkL19Wi6ssoF22yNLcnxioTZDqe0VTznezGc5lwhgtWGc8FRUvJS6
rdEWlbda7nsbX/KW+Aj5RmBqY3YVPySnrW9giwW9c810qX0LQUnLLdnhrD/wY/p8
ySmIYLek1Nl6VEgZvYO2XRgcpk9x+m2NMZaPWTJuaiGqnZPtC5gCO/arM3p+ASZx
Yg6S6JXfYswhcbhFlsHv79aea7hHbPn/drhhS5ov1mCL6BitYWwuvqhEDe47bro9
9hvZIHqo4UmB0XO1i1C0kT3RRUwn8OgOyGfOXLMQ8ptiqcxPpUckRe6+UCxSHIOQ
BOpmCv0lNETbQGGZzIUvoEX05faS0cRDyo9QUvx+SL/FIVqnQJZFk0l1wR8a22mg
dwmLYgbKFwJd6fh8xp9iSCAvJ3tL8wb49DgMqDUD/ggIR/MkZR/pdpO/gWXv9ACx
WkrV8SBj/G1DtrVDydtQaMA/834zyz85Gdp9cuICwADEzKRwPaVm+XgytJnDRYRZ
+Y6EpwN3AakDF8l9HR9jSAm9ZzWZWj/YmWKFnybsiuPHHtO+39Gynq4AnTflxcxa
wSaKfDw5quZPLmF2dcBEWb5bP5uPQgYu3rPSJCNzeT1P3Ic7h9Z1gjyxKYDUs7W5
S2glyxU8hcmd759eQ1q+f18B7O8JS62uGy5b9VpeM6kgM3P+8zX6RuynlfzU2IIf
BInuvkbAmDmi6gFsKWdmrinryTf7mYXqyBgtMAzRcVSAd0NCfV+DZX4+THQUIi4C
VH3ZMqYLJf0IDDQO7FVX+M763vT96rk1kpQpiKH2nnhYIYKp/Rw4vDZm210Lyul8
+iiweCR0iFnW13/of2TqKEAlvMJvN3coUp1xv7UWcgEXPocix+JaLgOOZBPpLY6k
U88YYTKrXAWKxbf9xZk+s/pediF6c0N9PUiQAiDrqV66RFrGCF4JQE9zED4j8gQ4
+07Gp8vR5BYyHfO/y5J8DWKkcaSUkzR8q8u0wfT5KiMbatNSrx2brUkPQq/4MuPa
IoC/XktzQhqafc6cqtLfJCZibNkOzjpNCdX4/VYyuu2UcYxeoE21c3/Y6kf2Lq7f
9LtrJbLu3ldjwS+mhQaBjS3Pnbnkv0//4A+enW5wjjOoS24zn9l77aXRS82ArGjA
2VEro66kNpoK08EXwug6iZ+OIvWRcDhnyYuWfs0nLHqMIoQu/ErEUAvLGp6bZ1xh
pxn924s92SN3jmzGxyk0h8cIKWA3nBLACp++o1XlR5A5u/lxYJAMrGA0s1kLyTZg
Kwi8w7tWsZP9WtPC2qee3psgJ6Ogyg2Tb6gJ+ZTGOZZm1cH4KtplTtNvaaThud9q
/Q/ZQ1iRkLAWSzKd9iwbuDUdbaOAgcC8jNvWfC+E8Vo=
`pragma protect end_protected
