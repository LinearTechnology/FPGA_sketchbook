// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Rd61Q1ihy4D3OS401KZuv99btsvubf17gSEb4GaHiRPlaGxeyo8X5a9xbU4qjsBM
gUryOjV+c9GsjUGoUrtTRx2HL/jr8nbl43eKFg/kbXMkKgvG6Ya+mWvPghjN8y8j
KcPJ8WCZhQal8VG74JIQIseQWJVAhQf6G82mlD4MEvo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4832)
KoNpN51Ly9wq2VE8x6gNj7mMU4jcWLEw/zlnA/hKK6TbGQqVCAI8pN7IOJm4hziy
/p5Rtsz2FKfoRnvcQeA3NHFIimMcJT4fmcF5DNUk5ZO8oD4f1p5YxFr27NUDr3T5
T2myE2cvx/Len7E878j3AP2sFr1/ivkAh3tuidXT459Fe7NhvaZM9SPBtcozX1ty
HFU31ryxCzi2gUeYRj9onBbTcZRsMBkAj6UDnfPkMOxwujl5v3phi9WUlnhPDnfk
SQSCT8IS627wJW/+Pf7rny2Tvom2JRQ1zXFIdZIoZ6oax7egp+Urf5At4QJeraDc
dbU0p4wiAUwGmJNSLuPf1K3YjDEW42Hr802EHtS/jV6BTmmuKrpfg3VAgZF0179m
aa2/wawnMj5sEd2OBPv1HQNkCRMx8fX5O/TcBeS5QhJI3MaBoZEfBdVt/0ph6Uta
Tp2/fq5FLEF0ac5Pc2q4fFVQMOgkhtsppwNuaJ5qjC7mX05/0nG+vJ7b9B9OjNS/
3JQkC+m2Zg9veo80v/B/4RWALwjyIMm5aVtcSx6mdvn1xDD76HtJtVNUc2x2oaSZ
sh5KVcH+2Wm8HTFdwsPeVwFI+RY8uwSe8dKBiz27EnuR8UHiYoMjkL9yzX6QrBLN
Rv4CE4nwdHEkVrYbVXig+iKHDTCUVp99vgPJs8J++NvXM5jVLWhAyDFzUUeCLfew
9e1ZznXJDmonyCGaqNvtrcjU7KSZBPo+UWgbYCh0ZsP6TqJfOP6ycBY2LV5M4hQJ
oSshyNO2ZUmyRmdib6yyzBGxgTK/MHRwELowbQ0qXb+UPxa5VaWgfgrRksnLfZI6
J+vq4/pY+zD2MvVX/L6GjqYRGKjDVAQOGIxCtxGfBp9K/DF+iU67qc8VuWRMAmdY
rRgVG6ivhCNe/Mk7ha/eBo8V1rMMYK1LZ2uWtOa3Mq5fpZ5+l2izsJS5WBkeCzOm
VEstz+0ymtVUoerkXdO2c1WAefhDHl8o6U7MHfFcz+MckKgElhEvrynHDcERjJuH
/So24dgRw9dWJMrEMYBvb0+jNQsIqoT7zXmu7LKy2JfUkt61ktdJW7IHv7ylFAr2
+gFj/s3RY52wETBeu9NF+gTqrJ/mnUyoDKXs8Z90oI8ep0dzOq2gK6SyqZT3rpha
vNciDQTJk1TnYUbmVAmksn08eZfskIen0YVp1qNESbrmPJSfgeX1tTjI4W0BTdVB
IYIOZLwElF0fHfuUBqXdpR2tuGaTfTzbSnV+tJyCpiKvGWtKwSrNtNpHd6AHH9Ie
AYyyqV4G61q44QS3Ob+smeNyqNIyLE7IcPfe/a8vnGQNDTmQjHpsSnDOLTf3odnA
4Nr/+V1H+F+bHO2xQsLpkdSN3AwYD7RVlyGQtHEblf7QWX7GKDJn8CiRbNXpL3A+
KFxpd7lPeugO10O3FARAptsDCrT9yLV+wGewB/SwDhYZ73arGuXUGyZTInVaAlV2
6mkqo0vyHKlR5vaQcKbvyq/lS97VlAJX7bVVPH/264DOqS3XrCmahlYUMR62ZcTm
ktxXiH/ZgaIrDgp24MImUfpho/Zvg3YsCA53QfjyYTO0X7Ed3O+KeL87ijgqFtYK
akEchYG119CwTXHMt6RIfF1w4GZlMtm3xjSm9f1hzRXGojq8k3iQEU42h6i+QcFw
0+q1wqWjtEs5Dsg5bMbowT7Aa6EfZ1ixNftGpL2WMH7MtpXXwJAsWLjZxbzf5wiq
yXcb8GzVbeYL6VWktK5lufxj46eB9nO0kDcmwYN5nXjmmiT0o8ISPNbZ69rZNwRU
DtImjKq00FlTdUNnckkj4ndgA2y9K1yrRAqulIaco/ACDXjfwtB0H8FwpZ1lNakn
P8zPKIdXiZNt7DFTXk31UVa94uv6vrNX1VNgORc1ntE6evUETBBnl7njS38u9gnA
s4n2AtgVO5+XuAgXk8V7mLwML849G+ypxtZzFM8YQRT76LJwnFd8Z1OqdVEfg8Id
huOS9CU04q3cydXJMUVMJf0SHSoJVlpFnBazL0stE7vU+yVByeR2h/W+JioOrZul
1K6RFJTtblfdlvpj/f1KXiHuE+2n2I7HLv8QlGFWKlBI6Jz4PbCk7UfKEMFGw7jD
507jXsiOHPD6DakhLAedUxc4VgEKgziXsLeFPxkl153cn5cGDbMvKJvQp+QR4gxB
pOMc2aVF01TNoIEvmtEBlBeFdv3PYlhTxscUt3aq0fQyboaDFWkKeOb6hy54kjVs
bBLEWQbv492VOD704F/7QVltERgYEW2XRwtrkHV0/sk5NeGhWahmIcWA5C32m2qw
if9myqtbVVGHqxOdjtboJh5l0YIDowT76PpXCzXHE88u7tW9KKlZj3KWmUfW9bne
/99b71kbgVUXHkx6rZeQKF1oP1uLxCQyQQMtsn+O4vMlkSBruzop2LXDdL4KBZn6
VEMzdC4cuTGkMnRlaMTtKh5ZfJoZp1U3vXxxQu1pfufnwJaNiQQ+d0w9Lao70CGs
b3rdMj3AbJdsqNFqQvQaEeaLLGWnU7p/x43+Yyt5/aHlbGAOuEuZ4Vr7Qj/M0cKR
j+zdNHcid54eZdD10a1CIVKV6i4878BoooQh/2eLJLVd81eD4ikABSq3qZ1BR7V1
zlPVOtGMV3aZXt/TN1uZwkX26AboFnlk+sEMLW29PIPiF43uhmzBGrDnXVjxUT2T
0mBvARYLaGfCiA4Iw87XCfUNM5gYBFJfV1qq2//nl5Eev72TuSf/zDi25t7fH8DN
w56kH2XPC79fVFzsqOoirTSj/NDWybTQsf3Q4XCaZUUbpOsjmX2Z5IFUZTuxRE/L
WzEUXDltdF1DpyIVNHD2vFQIWr0q53QrSYebPYlZAab6nBD4ev9kfCqN4Izpro4H
VdHndZWqQvkREqVvkkyRkzamNXH/+ap34xE71vfTO06abwOeg7YjdgWHKZWXbxak
pK4WeAwf51u7W/Hm1/qf63yKnERkvvChw28+NcLJvzbDBTYS7/+qBsZbPt0LrLvp
mBnVm1GXSpMQZTzcTxe+vROpscnFMxvoFpVX6tWNQvAQB6Oh2wfyWE7CT1ouTbxs
TnYWNszYb5lFxSNw5B7AXn8yAHA+waO8SI1HX6EuxmmeC3v1l7fh86fOBD+34nZN
UyD+I3XWtVRUYjAzqLVPCnpu7g4OnJf0slhrK9nC7CLch/pFgY+shw2Ch+dmPxsy
NnWTDg2wtiAIDtRf8WBkNUFemgGnnRULO6J5vqvQqipwx7v04qrbKhEOmBMsfDu0
yF+lVnHNBZvcq/VolPs9NlXgFK2Xs/ouKU3yNGYZpdL6EqVVgWO7/UeFRpOgkXNE
ZDj+hYWgq4yHvcZlQ+wiYjhA9iCy6ZhcA0Y5cy1N1UBhi7RqWBYdtKOm4EmI4xEL
NojUTVP8LE/xFB5aqO+jPlneNoN+PHfXUthDYNIAbcMYGBneAmzAn491SLfO1Hnq
TOXZi9PA7j2XC7tDf1rmf05dRJvmwEPa7rGhnscGjgpT8J3PmhMXlMZUsjtd1Cm0
39SbuClVJFWiEGd3yq5T3V/sft1p6y4444Wv4/sEQdU7hVe6LHWQvPFUgDnT+oR8
Zgr+0NbyRS+4PbcP9YI828+r4XUPbchPn1R28JMQMd0R09PB5BqqIdP7GJmLelGm
GQfH56NxVb5l5CUB1+0lsTEQJy/2fyGwVy/k1z/ViDvJBx7FoW6vkruCXPtXvC/r
ardOJxHsowvkUsrRelkjvR6unej18tWBALUht+/KJxzN/tyeddqREwRLQCHuVmNu
ElMFeQbUKsnQSSFNfLRCBq65+zKHJf3Iq3TLO43ZMizd9YnMDuwljS7M53RTcbLQ
+IcuPz1RUFmVg1oF0RWo8QSNClHiWkupIEBeP2HIQgf3HWgNk05gX022cfHOWdlk
wTp9YamtpYYa8PnjBR91WOtjJwwI4hJzR0Y+oEeEzcUfQob88K2p9tfqR/VEZWhL
Dy9WJEYgSq6X4Xmx7k1LfcVS1eI89ZsiCOjaRuYgN1hR17L9Y5AB9x7WRCxbolQo
ivvvyhvnbMUbDjSd7jNuvcA3k/cF154DKPLyUKgpMeiVGjvJrF7EcyOnhS+HDVVC
5n6U+xpP/zeamBJ8EZZDZJo+ByUrO0EIWX1K1z1n1Jb4wlU+WJRBVbSjCz/w4z4Q
pHwQ1AkbBKkfeZVpPl07FfaqmCkzJfaaNG3bp6WiXvLDa/t4lSOgEZ6aTdvYQMox
ZNNgUcZPd0oUmHF8XomJm/SaZBzekA8Oav95T1tYGqgiG6Hfh8HRFNSj2S+7UPUW
88hPojnvLv2XgvkR28jI4KzAIP4Ueyy8AETbYELrlG/x6lOgi/NUwzb8loztW7rd
oC4NQI9QoI4m2gVcqrALSYzSi/5a6azNnopbWBjQbFBBTQf3nNKrQ2HdwYfn5Ot0
gb/SwP6gZGL6TJ61KmZ4Hmzpyg+fyxuDRqa3hKw8384FPOmnlOGlmAzn7bJLgMfg
V/DJxj59uolEObLF7as1bf9+jLPGkAqpRzznXQaKTGw3KrahKpPbdLX+DKk65XIr
SRubzRwyhd45i8HgY4zV7PGs7+F4hEPjPTqFRLR67synaFDWO+64CMrzrFbq1BuP
GZZQM/dVLZt5i7Zce4IJTz3mrZ+vWH8Ae4hUAr6JEo0L6Wk0S/HZEb7KcOhFu+Do
2wFk4n+t8EqMqXr0mLfnfPFVDoL74FmKSf368GLOscdVTvakxyhcziPUQVDNU61Y
8Rx3HbVyNbexlbGQ2jUVu3b7LD3mHPF4Cms4Derf0h8M1DPs87++HeOraLVxnO3z
e7yfk8/HqvK8pkV9UPQKskw1tJDG0K2jEGx9g12jaNQM1nw5fw96JlHHG2wBg5RC
jTYVH9EJc/XoJTSMny1/PAHQnRnwJDdQGZivjdgwUUWp+a2Cz6yAuhIfem+HxLRZ
cTygoErsLAUK0ujzCw+51LnGLCRR23Q1QotPAA4uCyXtvUDn75Tnhs29VZ0Vov8X
abCGeCYAKV16nz+SGHthb6t066t3rsX6Ui9merROxP+Tpu9XF1E72meEtUqoed78
T6seH34hDMbPYhBAYo7NrDY+kXhHPKSI2bHjREU+Po/qG6Ve7zwL5Ptyzt+1vQKu
FQdLBsr8gOpDJHu5dROF94XE9U8ePJBcp1tpVH2TPAPF0wM7l3kb3g+PDJ4G/RcD
CPKMI9BYYaMs3CUDaw4bS43FVSBtnY+xmQXQTN7tpscVjyzkP8YqBZW4B3V+gcGO
aNVLxgxGQULGXcZi9J5ZicxxzgpsNn5nyG4IH/RuHpWJIotzobLcCaEWZtZLjDjs
rFNkWRBgMNaK8e+DnTB4lbNCFWT0K8E/RS9daH/1wIlXGDiRvk8V3czoz3pKixiv
bBeQJ9g20sLB0meIVu4FsmRdX8fAM6TYylgiW7VKVhXWVXkDrwntbqdmSjWdaJUd
5hzEGrbhiVyqOPWfNSEsCzzlTuiqVOoUeciEvgMR3V7oGZHkkBwuSjJdCXKemKRS
4HGVaoQkKluYM6aWjL5zSxg4ESEWWLKMYKRZc4ql8dM2SF626vR2FCAu9bdfSKXR
fDjgoBqXGafML3NQaN5Y9xrPFlSYKyRW4cYVmqupZ1SDxin5Ii/s1rYFk08dwJrK
MutlyzwTuWjLfLJCyzJkB5dDz9K4iwA1UqDQveBNyMiObOhAlyA124t1OG35zmS2
18Tgw+/v5jqG86vRuyXjyncKGzrVCUKgHzplwyeGnsiOTlABx9zCbzEEwecfFdqV
j95NZ2QhkY7TjEtbUH0HPa850n0MC7A14jcuWlvU+1HCHR54BN3dCpLs8Yc/Zwqh
Ra9Zsg3OVoSKPLfcVXG4jvSuVtAxBKnAst7NEvdPSWkLfhufiHqgK47TDo8iYNuo
bUqF7KAAfCJ8BAN4BNeELjPVUPKvo4VWfDlryJbs2mPhhLTSyWIAQxmWyuQPEGzR
5yJq9883GFMV2rGquBE19eK0LC1iLZmwx/KCvHwVyaRlGcYFQHppnEy5hOp1Ne8w
0NRRPoDTrrORSxKlDu28Ux9BGwqTQ39U13uem1oYXuCtQ4AlTo9lMlCUrSC9RC9O
qFV1oPV02gzkuyZchPg8cvpve3GSM8emBlqJGh+0tICu90hmw4H4nR6Lb91f1cV2
mRnj0oNeAPWViPojULPXaSozA9fpxzBEVvP/sMD5CjOo2RNgcqjzKWUiLsMy7H8O
rZUaji0fiSuL0hOFc0mkGhQ+Z9ItM4Sg5+Evb9bhffz5QgN1J14xZIIN0LWZNZEm
noUv291WPUR3jE9BMIPkGZ293FVtIgc9EIB4apbN6MShURa9+EGC0g0FbzOvnkUn
6RG22cTEYxhcdjhxuoT1SSM30TcxkwXOoImLFee5QgjI7zKuGlz5fFUoq4Q1wTEe
0to8f+xA8HQRc7XwFPj3Fg3d51n7/XevhbaQ/1Iacc8=
`pragma protect end_protected
