// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W4pVqzktESBsXl64D3CeiDA9w83QvVAAJiepQRavFQFMCCU392vgfU1XPJFoFWea
bOXaTtxeIbEaiklxhsfnQ74gEM+QdrycUXWRSLsW3ELyjXAzwM5SehSXWTlyg52i
GGEmn4t5ABZ9MFGc3FCen82NolDESH0xOw1JK+klY/c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70144)
Ei7y/P7afLaUP/Yw50FTBC0PoxeN/xXA9658KI5ZPuo6MIKir8oy78OD15ynP5fb
HlB6DXIr+vzNTNGRRtjzazy9q743ldCd+UIOXd5bdmSW8h8uKNm2tBpzL+h0wAHb
GbrcLGpmX2ojHqr+6RzoGkj3U6LJ5LgTuUDYxT0OzktH4+p0MWpoMtD3HfcY0fvH
U3hwuLqkyqLGBIPUWX8/aBePhsRJu+N4iegWQwm11zIQ20OK2v9ws5ykR6j1gvRv
8wi/dDMYWVLlkZ/K+7QdNmEFc3vr5/JYmX/MP6wUkURvS7KP0WpkeCM2nHh9SqOE
GhX7LYXHMu4QAgwyq8+OzZqieVoPEtmfHMGe5l/y3HQMM0pvYD2cyfId6/llXGjV
1OdRmi4RVL2cF8iwsoCb3gaQMIqi+WAzJ7qW8p3dShlyezsMIr4YbHvQtEwji6IX
sVmzvJtSvikWiuZ/Ebc1b4xetuJjP17vV1UoCD6Ko2Hmoa52iNNVZdBlh7Bki7GH
m0oTJ6KkueYobB47pIoCKPpHXv1FFmuZ8pbSh8fbKCsp7zRCeJi58/giywlEMvtM
W8GB9DfPkcQjvGsLiyfM8/43dUhuUIlhoHAqtgdiyB4bgrqxnjG3KUYBw0PFaFGn
A845Bgb4oQUxF8PSE7VHHnJBHYPk+Kg9OIyzYT5muhHWkzo/EG6JdE7vEkpce5ik
xkeuXIji1ZF7e5GP/NPKqBVNWCsRFK+TrH2KesfCSpNlka4j2SWRvFU78DHVgh+t
mbpwM3WWcNbSCNgz76mhtHEDlUL+WiF6RbAwfaKp1XzbOHF+j+gkFmjDPFHNgq0Y
PEU5ms/+M/6Uu22Lq5DPhIORSccn1XlN/sdaGcGW2qLHYbcCIN0G4miZLtwPCW4V
1gK3xg4nn4UB94dM4iU2WaJ2ZsOP5D0rc6LOCWPD8LZFgubKECU+Tp7A74I3Ycgy
EcgiE9klyVcEG/Ih/Y/9QQpdnSIsTdUG/OPy+9zDZMM7TKvlbduhn8JriBrBKhKW
4HsYLNVZykMrxevqIiTsXUfeznGdqFUtPFvxOiihmItGZ9s5tSaialFrdvEM4+8F
WHOdHb14dWniNpATDKH9AvQEw1RPCkikatBRfJ1dlbcBpyhQt8mXCiV4s5SnI7F8
70AeRCKYm/Hp1C81CzEWXbwS4Xh3Y390hxDKxy4bsu72jlu+BZOBvlWPjwcuY2t/
Mtx3QRUwNAOenMbhuzP9xIadgGtJNKezE1pBWOUxq7XVqNUY5bKvkYjQI62MB1b5
VTB8oSqQ5N86KdaX7cYa78E/knOzMiYBNfhwTeLA2vQ8d3EvGg0oc6GCeyNDUthQ
0vZfVzfk1lDfKZlQiU8qK1h42hmjPNZKI6Zn2pqve5ByLF3ladXzVO5apfC4J4YO
M+ih+Wi8mxspGRUMjwyaJil5l7RphptsM6sfKOccQ62qMYYskfAnG/dqbGjGEtxS
GeHrd/pvEl2plPPwlw87RXT0puZWV6S6Mg/V+nTYpAbhFSrN6EbmQO/txz1G90Xk
pQ7fo1V3uQAz+HEs4hkitpxxrLdr0ryy3BzPD5ZbF1/SL8UACpvtl38REJ1raiqK
Lt7aSj4dIndZoJHsmsk1yDmlaKrW/l/qDZ9OGccXkvjxuZCrXX17SmcmByx8JD7f
n18fQNGgkbZHVvizcEFRiTFKljXJlMm+3IxomTexDAyltCXE8qqvpzDH+yqRhuNq
7dYLQ7tRQ5/tXWRnReV7SMUIaQ/8WdOrop/gDkBqdocm/93FD3yu+dX/kMPXr6TN
vQaQrgA0DLERbXSj9RE6TT45DNX3CQK/Wku5v9ne8dX7YGzibZqCP2V3ioqVumer
3GLFx4DwXmswdP/FbYLQwo1d4CzyTOCU9SdPdGkPTUhGkgCJgglfijo92DgHTHRd
d3H18EGsHWl5I8jHASLpQeA4+cLRFgg+M5xby6eW5sKwf95cOBTAWOoEH/dUXCEp
SC7K4BkeW9PePG1fPpQCDTxVDTahjugD69gCZM+3ngqrxp9sWU/SwgJ8xanJDkBn
UCGFPNDu6JzEcyTGNio+piawli5QFkGPE3RDDKtGOVztvGPgzpCUOSN696RiVr7z
Uyu/sDdwDKLafJ/plouto4fcyMW+f8UIqJoEkst90NntoSsJ0+OuLdSldGIdmvfN
lh/PVXwBD9KlvG9pd5Y+AXLAKJpCPlJdEcBU52HheDCHigIGSdk+8HDpgpVt4HeM
O/wNddO1aRmd2Vfgny3tF6BA3HJaceLm/whfsnmWKWTRzV4NIqORy7KqoTk0DMR/
Is/ltybWqJLoMaPL+5h/3D4MVWsmNhbbvexBRuA9nrCPrsW5G0C0SoE3b0vutRON
qaBVr0MHnUVTzE/Wyhzhk4g/r4eA1B2fptKZ4Bz9oGOiRrSWPyv4L5rNbX3oZ/sw
uF3vD0lnfW/yKZkBNl9YMdoGd0JDVEtXyS6IaBjpWtGnptTJd/c+V05R/t5LDDkr
fUTf8aPMBP5UOlyslWVp5tbgiY7lspqnghUM3x2QuxmW5W9dar/RG5jTlqy+Ltsv
BrkjWEWyctgUhl/qlfRE82dx9o4uDBZ9Tm/of8XkP09aO4Sk2h00ItipCahfrXiU
retNDL5I2OTfHG+IQb1PXdHsy0zlTXeMm/W9VW/D1ADiM48yK1B3zXRVPqMDuu+N
eQp6iZYOqOsOFCd7JO0GNDtConzRoHIb0jAak+7m/Kbr2+nG344yt/eM3PgIkCvH
jFX+ZS/QljzzTffysbXIh7/RpcxuMVMhzGeHiwuHMYgdOXRt1RN69Bq9+fu1n/sv
VrdI5kG+x3y0RR18TBJ6QRh2BWd5nCQm5Ai2EtuMzyawsYCCe/1/skLPIpQDu2Cy
Vd2xX1rFf32nOGc168yzdl7IcnrXNgCkYF2pb6ZbdRRlC1jr1his55FzS6esdEW4
ojy1SwJHjoqZfAVGsF0vGaIwTIakElIigGfna3gRifnbZu54MZGCipoQD7zlHMoi
fGg/hziaoF4DbZ7Y64tZsC5vDtHoEzCASlxf/QeXeYvMpQmq21ABGIb5FbvWlU59
QoxmFh8s/4zRoX2OcBWRdwPkr6enPlUOSk7FVipQMz/Ov83YAlKyu0rgaCZnQ7fj
iUDPvbTwHlnbubKCnkVqGXAbWAaHYVu2zqfjxsogbO59RwZYD+Gw9WY6ZlVROCs5
J4KYGZBrrhD5jB+u7CSU4XGnh8rYTxbyHhR72Abda+T3/pAfa9sR+BraOVbnavp6
ovQObgWMDI/yUVbFu07NuxkJoeqKzCCXBT6okqZlMTBKvVGRNNwWmWxOimMzUuiA
wmczMhNpg0i5CjtUNtnyWneppq/CmmG0n5M4csYiQpw2zvjdw/QoaC3prwemoNYb
IBNyi7V3Isd6U5SGMxlSq0ArOBwJ1oszuu9wozrp1BPZg09icD3rvO6hgIsXAAHT
mskuV4FWKWHGUKc4B35YBvzL/LftkLOiIv2TFO5k0E2dDVclOIyX+L+/taHRl6Lv
JJRdVqrVYIhdRdzHDZHd9wnPJ47oQBiQa84gn5NL7PHaf8poRWC7fdxljSqLQHDd
qGBkMd0tlJ1GE9l88N9WMTAzPpAl5q7xrJrU3bi7ONtAVVxk2n19O7l+nvsxBZmJ
XfxgcugHq77YdNMTT3/FRmYmwT7Y1PczCuMPxSM9e0ig/qXhrRH1IAFM9LFuMo9D
s2bKSSACavn3bu8Fp9ASVQQy9JZq5l5U3AOIlnpmCuic52gGTnV7qfqRtdEexRKD
4IMuFWWuKk7karzT8rER/wpW99P3P3ETcjXkh3OKyzIhypCEfzyIroHZWUP1Rj/J
ly/YsEsgc3AZoiaDHJCQoCdQpjA4MCwS474jLtipuDmU9v5AQ5B2RqmbARXVXfsU
V+tS0oZnzC1yO6YU+qJo9zsmch0lnkdeO1AjQwiYyRRDEsioHtpXLK859hp0wCJ/
J/SJ4mFGhu3qZ1plcTIoApNmz18hxPgHw1TnaGfj3n8bdRfmmfVFRyVOAawMD5dS
k1rquIs4nxOtMEbe/k5/RbkYYnRNRdzb1IwMVaXwz+H8vuQYTDH7+VyAbSrOgDpq
CCtyQXTuuGr2ODMVc4hALrV4bk5noi8Oip1XkekMV+MgB+SpIj91FTn/Vvhbh8tN
KfsIs7pgp0Jo5+q/SMbF8vZoH9LJAYUusq373SvjHyEW21lgMMlPnESUZtLd8KjJ
Y5t/c2zh8Osk2McvAu4tOMr10Si9xWiT0QzaBRoK0HfXn6Nd5SOrocrwp5DWFdzS
7w2xnZHoSjZ7eAME7fAolP1gjQM25wAHsaPGGnouFs6VKp19b+ozydNWQc9U/c8a
GSshiG3jbjH4+hSjSvNw/CZ1r8Dh0HSHAbtwir0S8i6Z5bCQyhAAj0LFKjmaaD6m
EDTbQCn0zFkpat6roFtGa3EXf4SSmvH/Il4ZQpJdmZyCkJU8mo1+mck/0eNFd0fp
5A85QwdSEicqBQm1XrYLu8t08pTKYa8lvcKp/QSS+uTv8EtHGpQ3NvuzVsD8Jyec
hYi4uWlglokDh5OJHEJDIebo/MBr24Z6EpPKVmLGcj1RjHPqryk7lAah9jkfUiFR
/tmcRXyDSPySgiI3sSd8dZZ64/8YuNr6vABVS1CHUEds3/gGA+C9YciSPHtWXJgv
cYHJtv+PLViww4Zc3CZy+GxSfDxNApdZYM90+Ug+KGZBRClC9K7GwgsEf5O2CmTs
uhQ+dSDhak+p2qthQLdoQkz7EJMaXnqBWs8IQAwiIaetgd0DDHLkxc/aLailAy4R
I9yCzo3MlsVPaGTRdRWRPIHh2prVIjX9UFzqHSAywUdGGEqUKrclhiOYWNwSZVgA
CIMSJ1nCp6+EWsv2vgMPtzFlntOu+j4tJA0yDRti/TV8YYyz2jNC6jww9YFzsrgI
H1Ux/ajLzwt+S19a/42eiRagi6Y2mjZvnokTiUF+up2hmJTLhxgTMDjt5nXGTZTS
N/ucbH6unlNq3cR7efwR1YeH4QbFXjQCzvF7tIK9SPPl3UFXoUIf47k9Kh06FO2D
HTJAFQS0khko5MzeLXMwSQ8PQOXbmhayDvfOdLcCv25QsRyFBBSfNFIOSFJyCxDC
zoPHJmSCGDgb9fwp47tPmPcNjb3ruGl8W4wLwgNagvRDMa1KiyDi7NyZJ8xS8q2v
/iWinlvoMs9xMyyQRqwajZNxOZNWbN9xdPtMDaLMQoZkE2JAaZUjrdDSB/741cDw
CuRh12O76DYF5BPfayVQjasow0J9r/0Cz141ljS+e7vlyh33aqKY5ExFMkW17D5D
1hlpxee+IxKUg08IUe/CWARallQk6LuoGwr9W2cAvbHN/em421McGQ9z96vcrTD9
9DsUN+wm59/LYhAN4xqPIMZgMa2vLemWvkjYeGoNZrHk49MhZ8ttH+5nO9M28luP
C9qEcHuyepbasWo/e882KbnEYffBgr9kQF5so3VI51jxwUsscA57HPknLQp11M3B
bNVQslJll5MCSf0Xtn7zC2dqdfHVdwJAIIhz+yzyWPjC8pBKmuwz1oaTO+OSch/d
at1j2t0SiqXrMaVMC0/1ltRMFvIBdD+UvFMUmgUxDKiMCfStulizJPvClxBa0ZlO
GOxapgkX4z4ausU/emLZPNYBLGU5kFbXKJUT6HaGYklodVNYPaGjz/Sz8k+XAQa9
gr4goGX0yIPSko/nhO0J0wfJptZr/WpQym96cUMJ+hTvVvKrtyp2Av4bHYueEnHs
Sjh/GIjQCUHmy56Nq5tNWsZU75ovaOW5mJ7ACB21rqY6a+lesHoq/3F7PobshsGK
lMTB3HAX01oPrj7iEaew0ja7LDVQuB7tXLb52dAIUGQAOH6ix2DgeFt8aUAFQYU9
KU4xCuCpfUpkvXiix3bJ/ItcDhg2F0u/4e6IqNlBxqmIMMNL2aYNg89RqMS7JS+X
97Ca1XjYU4jY6lfRvcyvE3XhYCZurqpQqWwDCf5+c17R3yp1SwAWgGwKSIAo/5W2
8u+2vONEeUOBbQylcK9sAN4Z5s+R+4O7smawG1gUT5V8XI47HAr0G+WfPerfwqbc
omS6ySUGe/OTbBgaYxqzab27oBzUxzxIVl5jd6FsYbZ+PY//2A4MeySPfyAT+OP3
WvnEVCTHMzeLF6pX+8DazfSTE6+jYBkgZgJ9iumBrgtm6IF4NfjcydMU/TvpJnG8
kkimjOi+JfNdgo39yJ39MsjeBZzCci5xEwamYr8Vg97ckIhZACdgShLV3S0XMbdG
1TMGE7jSuGZsqu9B2e23FETqhjrR9/lfzbTDj2S8mf855e2FDrN0dmpsYGMvK+qj
UAsioIK1IMASR0St2ItME8WJ496V1NpDZrmuUvH3f/BYzbzan63gJeFsr/Q5k1FB
xSyuErcJsLXxw5OdZElfkDsTBotXFi3L032LEnXy01b4jCnIb/vE9mz1WERWibIO
dhEE4ceCx9AECjvJC/bEJm/Agtw4vT9SVE79plmcLmq24VzRNWWxzK+rGTk6Lzhg
R4rIt6yz0021j/THIVLv5NNMNprKkL0BrG0dRQJ4w/be7jHfN8UFJ5UPI7aL7oE3
cNxmTSJ85wdP4NfX0EporGw3ykilGk/Lm8yaS98E/iCrNuojuARoIpOx53b/2E7w
rfWEidMwCAvq36UeoVZ/O9EaInfg2BwZlUU05hm8yXpAhd09PPY/cWfZ4ZriaJI9
NwpNNcNCstmET5vF20apZV/qaKfTGQVD29pl1+RCISWcqfE0EhNJNtsmTZ2Q6ssd
ODt85NWUlmvUnUPDe1Cveq2YIKPbK/pE64HVyHPzf/L0LlY61KF3bHoJh8mlAuTF
J3j0ba4+qpENm22FY4opt7t49eicD/jxJJ7CtGCiE5CjHsIQbZy8yoIu503lhtWk
ouboOAxlC+7OmDrNIW6I9DDGeTW4/sQmIsueEYmRH7Z6WNfqRNqxlS44oN0Ma7gu
s6CSq5QKEIBc4ktnXhCopFtrTfAG62IXI8bbuahpQFwcwElPwzNu32AQmVqK2epr
K2hC3EgtYlQIxJQBVyaBuJOq91HVqj5Yp0Lfy/fgSUP1GkcDikpU1mQVj7gGNqGL
xmWNKdSzOvDldSIZ6+3g1noqr8DQNBppHnMr1me6j2NBWM7KXEQ1tOe1K3L1ht5S
EQ9iq6mMa1CNculwxsLcDwxHwEdJpYQxtmxb4V36OgNrLTNlQr15Ej5QD3a6K9tt
H7Dq5yyb/d/ISG5hj/171mI/+uuXEiIJd+Dtptl2m7jrTrlcJxnSCluShmOEH9eV
RrpO4mdzAwxDtEtifucDd6JBzTGLxTUIS1iHXkRjByUAIpROu4IS1MHb2R1NzSFf
9XXPUpQMnKuXFqCUsynaRqlCOXp5ge3LMc4QYTI5MywMIRrJyH66+1RodreWNU1I
IAK2jRVRZljFUOjePo7KRUvfxXtb6gU9QeqFBiaY7onKp25w4D8rP9DT7UTTwvps
4H400WPFyXvIPr5TqJT/N57egPfTe0J5kgAJalUMLXM50B2X7cbv3XKqdnmzbxaL
wqPNOwvtYrKgW8gJVVmmdCoj2oYQ95+jSAtJK+wLMMMM6yiHcbqsSJ3jOEICS7c2
6jkC9ZJpxK+HDoFI0z8+CGzKLwJT43plywXAlGirXafpSdeMzUEjxnXnuPeGBlir
8zPjuYnihxe9BdqiCkuL+ifv1UK3OWVwHwjf1AGN5Nx/soT1Mmzi0fqs/gzdSetn
4S6Ge96E3c87fj4qL4zOBUHdvbpAbdtqiZjAAIT4zwjpBEyMr3fI9xJd3H6WFls4
QeqhxIHb/Dabl4hmna3EP3Xy739j6HKq/cxtus2s6LHIn0Vr1LFYfQn6Re3THu2E
CsdNqqmA5bgxSG+3SdZ7dbk4kbWCcsd9lFLo/lLpujtldZs3ft3HuheYytoDj+96
VFZ7GfDIH9LBQoAZtk309LwNw9utdJ1VJ3ohZ2SWyVpAwSax65wmhX20MuYgpDHF
OHkMtsJz8R2VaLepgstRBXFf+P1wVa2Y6DWFS1grQxR2AQfZwmmD+sXZl+3GNECE
roqEgkYzELaKxRTlxHlOVo2sgDolEf5o/NhuJZjAY4+xaEaMH89uYWdGX5pMb7pm
Y5oOQABZ0D/hqbmrswjyRU0oDaDK+mcTwSqB444p2nVCGl7/vXs3NcHAwRSNxo1U
GHX7e6uh2u5PZavqCsl18Lrqzswh4qmR0WszJbIVEleep+pyH0fs4k6ctlI34RXw
Ul7JtFfYCPu3/r/oGuGXFjbigFjtijkVaF/1Z+yP9vf30b+giDvax73/FRLwVRDq
UWIVLXhHfUIfQbBx5+NUdF1dTQKIXQ7PXTm3Z/ZvuJxSADRJWhEE+0zaMR0ubqAP
DkMkD61q2bNkLkxSGWjNc1wqFgNBUxNwXpDIInl9++NtK8WdDwwCaDDi83fufdF6
NKuYytnXoZgHQTufpo4tNROfBbh+4SC85QT9JkkoDJqGpIZ+5Qb6OSjgBU6vKXZk
pzsZ+rj9SsDCM0weMRyxwsG4SHoEx0j0WLgZDRd283K59VkMclqqVhUyZJsuoLzc
xHl2uhQlGZv5vZf5OlXEC/agnHg8kLUazFCEdeJbBm4UU7ef3IuI60J4hsgG/TC6
vNGgju+RRFzMHYnxB7lTzVOsQhKXh6RDMn2R6ALhGQZnGvtkJBLzVtE9xYKsJIhg
5bjprAbSM4bN/Xbx+F/MmZmUYIOcnCLb34WAwROw1wXYhyEFkkv1vAuj2vkx8a7t
Y20eRgaqtlf5Ouizbnz4KAtQN22vduD0iDZoXe62bar8lFSkI4iQrfRjz2FqbkoX
IRv/GZYnnMgwlwe9TDGrbjXWCVcJVBLZOZMXxGbAv6VNPChISbua9KFBxECle7cx
4BIp7VEWgPEbZTMgeoWbVqyRBc8Z7bjpg9rx7yvClwLxgodeqTlH6+Btq4UOj4YG
IxX8kdzO3zYaZ0GnxK0/ea7UiNhPI/j9p8gyQlgRPqMo9Ilb3YYxb8lJbsMlxP5I
aX0g1miKKvCNVeQ27TUmiTle1QPDHxJglSYc+aamf4wWkZ/EXLtZEcXXFJZHTBN0
5jQzIYeXijJJm4NLhfND0TWAgQ7aynjys5mEFI9Tzc78LLgjtEqAZeAgq+qh0BOJ
cNc4czsLxIKMZxJbfjUVJCm/WhZFn5tjFvpkGHKTm59yTVbkOgQq6PMRVD7C57rp
WPeNmg7ayB5o1tyTuecMFD9jGN6F2Cftvg2YudMBAEMwt8vdmy6aipMkblKPh0ef
N6teI9sDqdwHvXcO8qhlIaXliOD8F72PWudDYGYkxPwZc5i8CkVjy/7YDu+s+G6Q
u9nhyMsM75ouQaMAnYqUM1OoBoPQ6JabRHG/njzYGuvxf9u4Sd6SkbhXPZtLEUaG
35vZEZpqkT9RSfL9vMH7oHpDJtZzHdiue/K8iGy3vD26aNmFdQX7FOToX/mYW+re
5AyQKQVaVwYnwbANCzF78JJNn36OZVk1NtQ6RoxU9UNxK+NVNr8uxcItpxj9+1PR
bjhX2o3MviL1HBMMWoc3GEsD2x57dvRAxHq7GqXDOlQYmhpB2BX89UzTqrKi2UOY
uQXGJ3pQoKqSiR64oG3m7kEluo7lHsoku43NTa1cER75dfvLWJnweUsK+suWITk/
V0Kl8vjfwMBGzrozA29Y63Tc1xlpbimX1/P4EtIGkrgR3STYfdY192TZKffPf5+U
MTR5sEGH4a8M6SEAL7LFJ/JhC91ryEimlMD5aF02CkjGTHznKGenNCBi/DZ1q/4N
DrlLbKdzM+VNHvVWZzq7URGvAzud77y9uUwMIUwPKMhv2tGqiljccmztbNYJqNn0
2Ae7oB1FydsWl2hSpcDieqnITcn2tIevAXaQS22eklTSgj0fiKgcJ/FGuHbHLBFj
v+Mo3xTzmSi6ZbbejCneeCOBKA4IPtQoeFngJBK67brWN9+fvDMf+9rgXCxn7kMY
r9SJTudjNNZ5n/wGIq+5uFiyshBrbUKSFfYcljQbeszANTlA4svFf6lxlPedyN97
0/BJmzqxG+sS5n07wz53cevRYYQrMhJh32SG4T/1krl79eg3RyC8hDZYxwJDalK6
6hlBiOp1bVnt+n3dNeGXMSBdEhz9vNhixgBB3KuinFNyxgR1gM9Te3ZNE7/2hqCB
vUle6MIlvxPvREN/bO+I62gaj7ez97rw+LNyV/C9sAC9vD8+SrtJDtgzHnq6g/jF
MRhDp/5hsRqPAKpa5W9FnBh6Oe4bFQyqxyoxGraYP70zhyJKOejffak8ToVuCYt1
afG/cTvCPiLzNRh+k+wxxgHSQTwVMTOKqv/2X7+8bADilyxyFNQjRAHey11FiJbd
7uhoAAF/7Y4A2ZgRKfb/Ofp5yIKbM1ylH355a+zSOGt4Wo7UqDM6oBBPSKxVNBYj
hHjZuU9WC0Q1vVsITOl5OM01+4EwtR9063BeQAwL+k/XIkjiZdK4NRGOwVgjtaoX
MJuM20GK3AZTz1NmbgH0NgSqWWv0oljkgFDaUYRBScnfOW36nUIRmac6p/2XKkYd
4MmgJ9lHDBD8JRKt2pE9/qfxhp6qAuS8Yaszmh5q0wMV3+2ebRXFvYKcDsZoBAtm
AVy3jPfx1Jg4mfQN9ISwO+Zqi8hDRcMMDbV9vv9/xwCWPgpwXn4+TnJ9l0dntOnK
8MOLwGmSmbMTrwkZi4cGdT0gYsibl3IPmQJzExas/Tf1tPnhde6TTBHyh4ffU0gj
FqVztwTuWC/iekV7k+H6pTsFhJENIpkGrpafS7VQVLXeXNjN0wdYJQXX7OVMrBwq
XyPgtVxT2NypT1PD2wdraRGXyrzzTDDYj/u4k3t8e+8NoM1EqoJ9VEZ91f8G4VpY
MoZweYaZgbmjXa04a3BYYEk+kolD0iRH9Yqdv+T2ahqPwYimfLXuQBEcwKvLblSy
dcA//ZIfRxBN9u0AyHQ5dR2pSQVFjmjXdlrDKz2vni4M5DKreRFOQ3wFwBI/coI+
wX0qXct7cnubROxPkwwd2eDFJYUtjOIn+wepQfF5EC/xMnqq8kLsQ5vczvHR/7O3
dcjOtI0KTMx9KmibBr7FF+owFazQmiRfCDRsqpMAkbzxZSoSdbKpbIsbuHMnrR7u
C7T6sfgZc7BFB8JE3tuj8Yp3bmrgapFQnXwpY4io7roerZPBR1XYd31VN1Pr45YV
XMrqkO1M19pZT5gEj+OsRYR0yR2IR/bxnV+QO+9wapZaPjXTnp1uTEtNd2aOUrB0
iTTqiTBroqe9eAt7L4T7yCAUMJJkUwCj1gh3OxNsn1vIDV7tiFJ2bsIDhqA3xA4u
1QYPf4osQ1wiC1GUrzp98+GucqFYZeqWgqjZRv1XH8Uen1j5S+4HHR4Lz3+0yKdV
KFh06i/RrY/c/6Wx7RQpwvvHFF0o57GaczX4rtaU4CZtudL0akJ4P6POkT+DmJZX
F8M05enbyWBPAx6329sMWjwcW6uRFLY3SxMYCl2C9kpiCm7jZf3ik5/LKfkathR2
L6thKobPih9+EYuNhXIKx53JeRpNLhZzQVZC+w48klzenFN4xVOtUWY1WlrMg2lW
zy5OGdHDFBGruukpjrwDxB+mPGTFh0llQz4fOQNxbqwP1syqlZJ4Xer/VZdT31KX
qgbYZhA9TaKIjwo1gPPrCSmW3CAW5gaH8cR3Ngb+ivsjbxETAv13J081G1lAgaAj
LXyDl9CMOd9/GZgQ0SdthjPe+eFhmBfj6cGIHkbZKgxxyWye82ownFB3zPSDfnZm
znq+3qUkJu6pwKuzqETSTKIIxyZLtZujCAelht50dVH8cKFoaYtPj0GsUbyEIf8y
YWLcuUB2VxbnGmBzgNmKLedLZjx0YU3FPGkE7+BbqOwxZGH2VKWrTlJD+UXZ97pk
RS0IqKs5oP8fwYbB9exyEEc0LBX/a8IE8hYUEMpucQO9bvHtO910n+oElXLVy+l9
ZD2bClcmLSGF12zwVk7xu3TZJqCiPtxdDzzp1OYiIC4iy99biU0hW1so6BHs7NVG
eXvPu1CcHVlhZUcFG17ud6+wztsdF+tkXHyo9AhIkjp5QpU3C+NZIwLJsuP/fIo7
8fE7e0/Lv2bzw8oY2GNKh9ZYVt/2K4nx+z434bTRHJ/4z99mmNCt3zdv4cOCkqgO
/nvLdXc+oBnCWKrf8QwBrruBOj7bp+AgcW+h7KSkZCCQtVr0+3nx8NMjDEXeiUpB
BK7H4xJxtKDtJBD6oSBsJZntasrENuq9CRWc2d+Irtc8XnmDuTAnDv417trXXssU
i/7pYHM3BIgGgPKnHN8h85Ya3h3lKzevBtMWt5DC8ivrRtResrRb7LsMgRR1JI6z
nbHEm87gKJ0hjNgBKZtRlThcFBGfrTkfCeUHINneBxl6ClcSsA7bURL3kuzQ0SD3
95/Dx7G/01rmqTvY5Ytn2ddh9JBxXB1GhVAWO2lBTSkXybHgXoIuAXgxvw5u+uB+
x7tuhKw9JVKGATLm4CYMeQ7mouL+WUqi+mPqdnz1QTHxNpHDnR+dUCQMb/Dc4xCE
Y9/YoHJJwyrzZo/Hrz0vRd8O7h5D+OAfkx865mNmMu59GIAKxDpFaHEQDdm2BUG4
vIVXYXBGkpefkefMDUfuFEsWaOlOCa70WxGSXw8kcS2GFw+QkyGO4dpY7bjUtFzI
1TgWJf4g1PHcVAVxBriVicYYtt+qNQNWZpStJMtOQK/JWikE5QtIimC92+qQsFLh
eF8KSToFHFMwAFAJPKRnGEuASqC/4+TQi34enOcffa+yqRwrh4CT9U+1oa1p84mM
Nf5vpFXJz6xBmGxCH3lv5w5OcuSkNJwrfoiDoX8Sz11vLT8KhP+1V/hg8W3XlKH6
qOnFtlXnrWws2Vvp+DJlQkbXhRkyxSO5lsuwF023f8WNMdO6FK/NduGa0MzNi3EF
B0YLVCIA+ZRaJ7Y5kyzA5jb34g9OFeaqYLJrqrF7XcABrzfUgeZ8NV3ytevyMzCH
13oThpOkihf9J4t9ELEWNxTRrl1ggk63b8rordlTvwO8FPYgdlaF1S3XPPzkiiob
RgwYurU+aFPTPRJ1YR74ULarDNTWBwQdrj/EgwtOavkizsxcKvSy/u78a6D4wvGV
VwrR8zkojN0HVSZ9PYOIOaIi8Z66Vyr2ExBSho5aDBFkV32KDuKM95Tv1yRmiV/J
ebZJEr1nEJp4h6vU79yyt71rzwFnTkNDG0OZk+7GTbRNbfhOMw/d61xnhK9t6lmD
ebZwR8YheqtQvW1dvxPth1Dn9wrUyThddYrOt6ifoWZBwOaGEwlyv6SD5YYwH+4N
LggsS/CficNvRmhN5bSilGd8pc3UX5iYPVKpT3X/5DdygLaWkDif0SIYd07v6xL6
VWrXXQPIJAhd3slwGyIp5JDFbodbnfgUjRKaBiYBOQxjy8/tQfGUdNX5sJlhPwbZ
xUEmh8vSxQrYiqoEHiGVBb2OGA0qprueeMJ2yvwiuJv171gqsg37EeHmGXIfoo0m
0PsVjtP+XUu3vbZ5h6hThYF1RG9azatu+H9AmxtYb1Ut3/fNB9shWs/ZemBUWSkR
VpXCbb7yuCUUiAZfyFFN7Yl71ypdzGNWWO1J2di6UILBcllfmZ/u2KsBxYs21Oph
ntwfCJP4dTmieCl8UCd7mMAQhVZT0gSkF2urtJSCzwbm9LVr3sGREOscGId/BryI
zZxHMXzW8ijQxrAZsiMQCfc1mzd0E4W0H4a1q6//L1ES4Zmbp/V1YuAhke8zYoC/
L2JjZsgVMGvhYlcavhFsfeKvUQouPf4XV9yNzwMEXe/B5vvvEMPyfe6+fKnog9+E
EsJqTWBnhLGfD0LRgyjs1KUmH4v72znyq4OvDZAVvA1i4QSbTwFMlFBq1ydLgkoU
VFn4KUXXyI/ZPSenl1u28WQTh/2+P4WRJ0CoTlJrX+YylnOsCh6FwaUWvDN+p8iN
zditMSW0l4gHFawCP6bo47CWm4B2+EEh7Pxy9doYlept+hsnWiIesrxsUB7YEtdw
Stt4wOWke/dPqzlGZoh1Pz/iT64Sx4jwqJ6YRsw/AqNhdOrb64zPjTaCHLPFjuVu
yvVLHMSYPrTGIZvgU4YoOFVQG/ry6NU0mKyJOC+PVYCIhEBCjt9/IAISB3+t3SM2
N37+74mqOrVQzs9NX7H71bw7owF5Dx/bL1jj2I3QcuJ1Jvg7mUgZDu+T+HNljnHo
aYwT/wI9m1vYUB9iHxvuji2GLoblNQpTkpVXo9j2ZnAYSlqBJNC64Djf4Db/fgcz
Nw59W65H950vWuRlJ+a5Vw5bAPoXIyETdRw6Tn/F8amceVvyLJM8VVpiZCSARa8G
eA31FiYoEO3Q7zVMmH3b+hkvji1K71W5owFgQ2n0RFMQRNAEXW5XIQp4fq9nLG/I
sF7hLVJ34EMMGqNEytxorV/Mqj8hO5jiGcEmymfzDedAA9Xt9TJcvbrrHtOy/kpT
hSwQGY+RTEbPG1juX+/tbKYnRbzM6bmGyDO64hKPUwGLR9Sdm1l3h1xJLE8kdDYa
5nNC+MS04W/shQWMZ1liKwJeh23mdxp84/u5MWPVPQfZZ4wA4HawAjcQhQwWdm5y
Z1LU8Ipu8xT3YpUD8iovGswD5UsK1oKlVCK3jidyhnv0RhW2u4cJwz57SJkwFXQJ
HD2a42D1EuZ71gXybAFFpi4xI2n5LHtE5y/J0LTc7N+BGcLhOcnE0XxhNCejksLn
wqubWpS1NF9GIuVWm0sVfNUj21tTAh1rvUqPJsn0fTaCoJ6RHHYJdD3MI/ODLop+
8jJNktKXeNXSBviowAQVqjpZwo0w0yBgLI1RgA7Gr+LZgXv89yUuQlrSmlVwRuAK
ECYSuQrmOKkd3V15cNwzW8UR1HyuxJ6RqQDUpndA7BgifWAK0ZEkPMp4z0kWCqPU
mbyERfUYP6c5WdkUNlkuKbDNHO+ihckXgz2abLn1J5irY3ZwRZ6L9PoSXPGPGq8u
EgCUECdGq8ZcQN9XY+KCn4aMobq5rWIijSrW0wqKSZHVc1SMqocpwh5oCxsERwJk
Ry5w7Sd0Y5NImt6zPVjpI3aKuXuOllUNPP0+lu7fR7JhqosaKNiPnO4vHtbWAmvX
VvubPJiuKj1NuTVDOdyBqknUtjKu3alzhzYj7Edm3Cw7FP5HcYBElH+Sgkbysh6j
7Qa3nE+tk5aCN/iq5wFFDGwD5eWQxbsYaA1mopqVbmjRz3UkeZikIyqcUJEB8IJd
lxjA52tWWac5EKO+sKrmgXlgTN11E81myTpeyY8I+ZM2RClm2lrH7fU+DjvKCMSi
+vFLRMpDfUnGy0STXrEwkE7voLLCKTmG/G71dMNW8KjhpU5QwWtHGr4N76/6LfnP
vkYp6KXDwyJ33zml8omD6ows+GhnYZSRy5PoJlYK8u77UbyOII4z6jX68fLOGnkS
fnQI05XDI37BKZgu4S4QfGPAqrvb8vcFkYpc4x2D1IZnx/aK7hJLaOfADOoSIKMV
v5sVyvblcp3rPtsYmnWG/NL0p8fDBQ9Z3ScbMABGWWC1euyNAeuIK/rn+U8BdeDS
QeXwWRmwb5BAGLmMerj7L4DwgI9W1fCufzt249hmOD1yVfLYiQmrXlm+qjOZ7Wfq
RXh+JEUCYzzYvfcbv0A6Lbsz6BJBorJY9Uxegl+NBFQDE3AoMLIf9NPJIDrvEtmA
bDh/RGDS6xMO77tzOzoqI4a/MAIvhRH/5IMpCj9Y4S0lfua0jqr96lQ0RO4yqRac
aJaNIBg5GQcV5M7v6lM/Yrf2Q3M35SZWNAAO0xyq3QV51I5dZOqjKOoM7SGSFCo/
hlETG3Hmj+/0WNqskwIqtFD5SmTRlfpTMiE/7jTmKm0Z1KgTHn6nOYFMaH3EYLDY
6F+60Ylin0w8woNR4WIUj8GyoFOb0L4kRQNnhowEk6GvQrUxhN5KRSqSHgja1z0L
cYmVE1CiGGb+S9qmYxkOkXCRF/rdwUP9UNMY6cQvqeP2bneTBjQ4m1V6GCOjRPTN
ZtkW5bT14tdGSIPSFmyUdlvxiJE4ZO/GJXdmOjKU5XLDQ9EjJHcHvKNOZqEj1txc
lykaARY7CrgwYNlL5Vl2jUgPX15681I6GUXEon0G8OEhoSQNpeU7VLnk80B9b2Pl
a5ZThSNt9QGa/YQGbrjX2U0+qGj6jEfeebHhqDGyyNf/QAjU4na/q1h+zkVwLSBD
lXQ/xwvx6kjygP+62EW5ZeuN9dNQ8yGgVnfKiiMCQa3/uRUfOLJQtB/H1+ZhDVF7
/Y1eQIs50+LKsJKtGqWO+ymA/3W9/w91ESzZ/zYf+XTKPScSxex5Z1PVLCo5rVs2
4Usrcu3HmQoaXN4M6reB680zdq1eedkeVAbKdUvMXl5uvnZ6Bv1RtFZq489yxaOm
9VCErZD8Us6SL7M1LxsPNqmWF5R6ezzW8WLVycSGUUHIzB2pWeM1NVlyeTp7+1Yx
r3uwGpDReaMCneYA7Q1CcCDuaj2PzfXOInYRFW7Uc8EbJrhHFDW1KCmg/ShduafX
wOKGC5CTP1afsFwGDPgIfbuLfR9Y081+LJWB/otVJVGBzGy1P+575zEGyVwgo7TA
756Y8U4LESTv6bsHohCQTv4e0SjqocaHPbGKua4bhHG35rfk1CAf2Wb6DHXF/975
HaZ5UOIh8I2RbgVcgRCVQhuYUcN4ivVcAme93um/3ltS9+SShVtpTASDFOlZPzJA
H7tkRSlS+wRwu+GBCdAqyog62ycG/Ca7TDu1Batai5me06vq/FZXoDGLE9nHayVN
PjzCW5yiLg5sC8V3B351YzcrZfPmCYLey/9CqrxSByhSqyWM+BtRbyHJyfcqB3Sn
pVh7u4qjnqKcT0Yo0ubE05vgE8D6hfPnbpRmqFIASpVSBn2CPuwjpqlZgprqNIL2
5wZBRiW0iN9TF71jgag7hcEYzPKnxae86ekKjn7PBA647q7a+qWAH8V5GOv95PXq
vePtC+orbNTbDotWzxhVyfVsOZfnjVESC/3Toylf+1auD5eCwro620aT/E6nw9wS
2qc4JPLvQFdzkDsGKlQkuCQbSf2p7pUubVNsbvGC7xcaiqc60or3c71zBA3JXAVr
SDeyPnjvaJjGX6pWntw3Y8LUCJO50bfHKa4EmPdS+zIHlw2nb8DQQMVEdJv68eFF
0EQnpzuxBX5FfDmT6j823tIzQHwlJdq0SYwXQCsNGSLRAmAJmCfKcVfG6Jz5wkSV
q/rGvpXHDWhgMye/c+ibbAtcOdMVAbiaMe8IgGG2bjyC7zkkMq5WLZSFE6hKArje
v8gziGy0aeq/A0aEnxZXrlKL/7MdG6+PA9k1h9QMiwRW7Cn3EXqdzCDkTJJl0Ctk
kSf09kAwC6gBKdydqaF931NuqoSBK3dCbsOBbH63L9E63AkbbWQzZ+GPELi+bWNz
FMFUsyHHbmC8JmBD/ZBRYLm9x0jIk4Mf2CYknzObUxdy6A/2WYjZBE1a2Si+WOfA
amF7glBmaYU11dxsCNFbxEd/GhAvtoucEnNrgV0pzvRWjQMgG+Umvhfr13bGlzu3
bREk7xnO2kb0jOqKzAtE4KelH6tWiJYdUzi1QAB5YZOK+SUVd779RcKEtTIb+3k5
blEDgbXUYONTelQQUYvJBVh/r9fxyjEuGVrs7EYpjbwp/PKyEQlv7y+T8p/P6Byx
/cvyipsboAsmrF51Yh834quvud2QRfLsC633zhkw8OV7pMsAryc4WDZyY31p1f5m
Z49r+aqunt8XQzPLGEWsrPDZG6wI5+yMU3mJpwM4hA8wGxqUsonmoRoHpRqX+OIu
LG3FoYVF1j8Djv8cZI6hG4QeRXjRbQ6wqJNJifFEc4dbjb0nE6VTEJ0BTNLIplRr
rHn9Nor+SpFA1j6eZ2MBuQNuxG6mjZbs2PtVPXybMMQlMdd0rvSnNVOyGpQVjexj
RIpEgxMJeJ0uCW9V6s7wifnRa8YIXxOGgqV8nbrZvsJKA6ERtsjnfOUq4vdxJlg1
goLuMN5PWk3lAR/8e5UXmKdBz0imon934pwkx5vSoTSqbjr8imJ2b5Ok69RAyZ7O
iWW0BLveKZWt+tF9eFxoOlkHeh+4W7xztJTy5TF9asZofkY5x7iwhb3Zw+7Xehv8
vSiRmLyU0HYttmlen+uHE5De6xB0G3Tt5qa4uPhY2azOW6w9A88vB9oRfkv21APD
2/r9He4IIgEp3JLzanUt+1Dj5IOvxrHChxudFDR5MolZcy2HjiUKlW6573ijnFJo
Mtfig3YIO23c0IbyjTxpEktoRP6AK2SkS94W/0y3s9vxIp3QyjvuA5uRspPho5kL
56GQAgMm42+OI0GyaKxxbn+FxSZ/zSO/rT4lVhw4oCT/4/TdBN7hiC+eMMZDpXLj
mkjdC3KR1Xpk2+OxMjI+Cw74W1+4vpnvQA+svDl2QJ78zKv5CdBrlOjmXC/jEVZP
gwLfr3WfO72Dkrr/RqZFJwQxgD3ze8s4u4bnkU97iZ0u8q+HHwfBofdrdN17XrGa
GgUjDg3dG7Xhbqli7hdB3cd4DZI6LOpdgqWcbix5F+uW6nxFBBiORge1BZSqAfUb
xkDzpxtMq4QNHegnBeVR5VqZ7KH8kxJWPnctug7cUX/WUnB37NoRRpwjA/4G4HUl
4GUvi/zBWGQeVwBxbAuycBVNb68er022LOLNAcL3ycmT1SY+LpTMTEdFkbaUCeCz
qh2yf81OR8rr36wiw7EnWdUThlR/odrxxHnMPpdLD1iv6mwQFk/Lvk4aJjFFeeXW
+2MIt2f43LyySqpp/bUIJb+tCpkoHuTPSS7BFoAxbPJAZJ5cVddrX0rEiNz/9r2G
KmtA8vCmuYEW0WTSNZt8FJiJjlCvEc+8wnBKEkGwps7D5JVwcVCifNn6b8i3Gbt1
jlI/+P2Jmuvpq/p6nUsKE6d1Sn26XUTiNqqQUQVCBk6jFbF28j0aKJ6EsrVE1+Yj
bFJMNvK5SGuKfDhRjs3t1VRbfzxlSQUffTksxqVoOJ4WhAkK7NPdXAFcMeZ82+In
Uhxi929aCQAJX0PyVOP4SC2M5r+HtMBu3AVfDh0MXA7T9bxJD6G7J81bgsRcIXb7
JOgN/UA62iIlBjh7fpQQpID19DXP+lBtSxJgIksO/wWib69wU6C/OI0aDYs2ia22
1NA0hTo6yf3gXkL4zZ2E/+SjtZ78wQoXLDVLZe0wW5xOiutNwD5B8a/p8f7qkc31
2moWwx1iaChkMANl+zqOa9SGodnzJTijtlmZ1/CFAkbDiMzNFjcAiahlgMlryRq7
IKJDRnuNeResAcYG416FZ0JX0+taD4HUklWXEF0gk528Xq3t7YptY6/WovhPD9dx
sybxeFTpsL4MRZdgGhx41QNj6PATt7bOoLB5nhrdh7TY73NKipboJPPAfrnw4qit
jTko9LzcLC/aibGVcrvnXSqp6+R1pt9z+xB/t+kNCjUDDTzv1YILfBnQ7ApTLbNg
2/Ibzpe+VUez3iEy9AdiNME//9wz/nek/FTNzl4YuwfMWChv1C8CDHNbkb1k9eBw
LQcqWKElqlnInW33HMykn9oqT+8JsG4yx0iuE7hcf7psxySqj9dkxQHy9UwoJnIG
z+HtU06QiPCLsM5K763gTZ6H0elu13C96/OoyrNzSC04iDNPGPwiHue9mmPwmtXN
QPcn1kvJkTWNDFOnhrc7myqDfU2IKWLu3Yeok8Tqmw9gUyktFmACriUs0Q6eAO0V
9pwKpIYyXiYLG7oB53KBsl2/grhS9hHDL+hLxQTq8rsh8ZhE9AwKfFWGctrDkuWo
dd7dnyOCv0RbJUTETAAyVHiT8XEFKPVWvp/9+n9/qjSxk+3j+CsUVLYTbO7MekjZ
71WxSJ6LwhQYj+BmC/6RADdESN4akST5WVBgNHdJ8kGbzp1ynvhK0IZMF/Lhq3O8
z2myQmfTYyxPY2TAjfi5Uy2Mu8z14AxK0CvHrjOIxOP+ugGm58FC3VtsGFnnz2vq
aiL7UbUaRut5O1HkrxGwrQwTLqI0NKIhdS9k1Nxt06BD9eEmCEnNuskArkcLS4iD
5Y2PLRep9ZxE6rguH0i3d60VBanwWfNi2gk2pGDFCvvnGUhSbtAzvwdTEdwi7rkL
TKChlhLs7B9Zrp3jVi2XY4njDi4aLab5TlcRJ6iHsotrJvMbrfU6Eo2YUUdUpaiG
2sCeIqOAccSy/PxnSh1VcD8UKyNoJIHn7GBy8SFTlzDdZEvkLp3E6jJIeNLqy+2L
OBw4inlfmQRJlKbCpK5YR8ANmpS5e7S/ZpQpDb15jYonPMhEIHnMoVcl+JihQmR/
kCAscgl8xnsDS3QL1hPuRr2VzC1T+vOPve+D+4BKbTQbqsuP8OmdyuoEQne4Yw5m
gbwqxrfzqzAcH7ZffQSzyf6I+6WQR/8yUfj9v4nNnRtVkNKD95uQFvgqEP0sI8/i
1AhTXfp8n7/gPTbY+trTAs1HN+pC5FhuiZiKoTKNCEMukm1VkCtjtONisrS4XXTD
mRgfBxukLmagLPIPIRZPDEBehqMRhDnVgEXVwRyRrKD4obFZRxSpoR9c+i1CQFv/
g8XdRt04dEBxHf2ThsrcPwGbvuMLWrrifutstiDSOlc+NHhOuvCWRVG8r3A8JY9N
k6ZB2J786XVtq9PUuYIVj4101hjAP4NRq2yNV9dE3i+qJhMpNf4iD4QUGMFOP2fU
P9f+y84cRFBWXbBlMs9s8fRb/jPwml05XPqrCCUzDiEmEzw2KUEKAzMupOWSQqva
kFB9PnexJCAHwAoMjMzJaj/U4niDhdaL5mKDn9JvlxWksRRvC/3BH/JLSLKD48Um
RH4N7Dyw8ySZzi9mvbwY/B40ROaPqtHWUnm68cgUSk1oAvUAJS+UAt32oyt2I3WT
DeHFMTB+MLCMy5D+JFncsKcoDj2irourp857+DnGNYNHfRqNhx40Zg9U//y/87oo
1XVEz35BQur9z4Tm4/71XRsUI413mk512GpNGuupm9SyOgvUYlmPuQF5iFa3Kx8W
xRhdKqrJHEOR1LkGJgBA/z6ZoBYA29zqBpgV0cHarlo9qzDu0A6Y0KjM3mw2UXvU
aziPhmBRlT9ZiUkDQgeMXd/jxu5KWKQ9wSWz7TrhwSlh49gdBALsnZ/ITYZokM3m
5nrpehZrA2qdaU3gN4//VfuDIZ6opWiDXRDSsMPXgaXqeRekx7e2pccQUzAXgP81
mp5ShGAC53u7zNyTXSc7I9Mx34xZh5UYIEkYF5MMeDkqjgkZXe9HJq1qxsaydojx
zejwhG9eiHrrw5g8c2kQl9uhaYZhvS56BZJsxpM/KKFi0cQ4l1kOcKUvaitcddEU
5X7l6ZInWqCJCjAgbH/RqJEfzNRuy/HydaRQXnqKKwlHbtFulq4R6moumpv+mqFG
z0Wv6MSUjyC0fwq7lYYmonRFXj7ayqeWBN8cWk2rvvWCmsCRfC1g7BpJgaNek/sq
WLO1iw+728dA/arfxkgykZIoe/xMNTpaIQG+L2HeyV3jsnfpSq1XETrXVGZAFWju
D8VPj2Gbkgmv8oT6SJ+KopxMA275ifbNeAET+YrItUC/DNxapvjOTffV8Zr8c3N7
2fBvegU9IeFAiPgfJyRfkfn+yea8UPRyIQrB8Ujfa8OpBgdmvE6dNlZZMf3NLWgy
y5pJcBhADFrj8V8ItnwBhNZZDxa2RrBr/qbHP7AoAY14S8hvnBSkqsqOVF0hvyOZ
YKJ7Ly6TKne1DKQkJBi3xiH9TbxIRTAgj8ADFEbDxF0inn4Fi6unkeYfeHH7LX87
4v2Lo7cG7EnEx4i6G4f2QCYxIuAgs10Kc7O8aYI/NIVcNd0qTnUy7PTlETESbay5
hik1KYqlKvTw58BqQ4lr9Ev17w+nn6pdxSu8gCVMz3laTLk+RERDtz/I/NSrAVqL
oeaBjrQY+F7ZD2tqFWvUBuTW1H10dy8aPyZb2jxzLKc7p3D/kbdUgQIdfCAkRq1l
bDrIrTmrRmYyBPwnmT0lklvMV9SQXLYm2sb/q0CkAb2segmRQV5CoPe6mIfOw1LX
iDaaXXAuRTAXad5/sdmcw5GHpy6DELGFB6toz2eJ0qHFFgExnsrwSkueILkG8O1c
/krxg7x3+18PGNfl0H6tqKTwpCofFDYK9tIq/QgI11lYRSLuYP6voUKjakzEJrnW
FRsDa9zaXSwClmKXknusdXMfWWEshSaWLtyLsp8sMUUtUCaMD5Tes2xxlBLAjgmv
Xu80KV6uIjxX/5JvFbVPfRc6WEbjfkFu8Jwb+L3lnpUENXYWA5xdOy+r4di4Vo39
qtlnaRIGsvgDoE+7glThosd/PrTpczxRp4YK5FiQCMRUIhi0jPhIY9SsyNr9nBz8
E5xXDgYuB/7jLKeVMV/PHNiZ4mhNiszNZwwfYRv2nQF9PRtE24Zsuo62fgNdpyT2
dmrdbpFp2m7l2BYOYA7yPUeqI5b7nVtuHpo6Dp3+oO0BtkNSZHOzsQ1Gx+orehSr
m02AY1XvvsMCwkjk7bsIc8jExEZ1lVGChPNVuC1LCE4C+0U08RUwTOQEYlmFSYy/
kASu5rDmoh2e4EfZbM9le1t0SYr7x2kdlfB0tMflP6e04ih/WAQYQY/vkg62p2rK
yC8D8rP+Gi0DUhNO3enwsse9dsci+Flhg4wyGAF+xYSXB6yNnrQRWQ0UNcziotPl
oH5xBOJEiwDKTdAWvQ8BdFUZ9PWjQuj3xNLB2UnApkEn1OYjb5iZCNto0arqCkDo
l05tswDz0SW4VCFVEENzOjEx781KDNVhiiXSOmzZVpcSzOuvb+Rfz9cupCsU5Bgm
25WgMD/ikK6XiUErlEgzK8IUTduVEEc76kTJzMPt6RmVNIasUTRXsKLX/Jc+ImzL
n6T9eBbtReAMxdW+qPn2hTSD0xbiWwLm6ag/bboVaDWoxIAFW3eJ/DWfKyRbrzd4
iAZZvIO/XUi89mp1gCLGZ6SqYens2GnQmaVCumY+o0eAM3vsDiP3gcLbDmGnb1tg
D/+a/TiCksuxJzyOOck/PFpQJJHNmsY+46V8tiyzLk1IBEKQTYDZPC8Kvul7o8F8
Dnh+VdRxi7hwpmSLncAz7hLy1OYUQs4/f/TffDTcNCKrdwY8iKh3pSXDPbfkylEq
juba26Hln4TmlusHk2q8CI2rNoWg5iSYKZ1x4MLoeD64iT2ThhpVnZ2Lj4j2xJ7H
CuooMnJNWQ0eFTQGTw04mWoTsjyDxoBDAWCtFbu/73g3hWoP4g0WNwf9v/2vo5ht
2Bs/YiXsXUPfFgEAIvKipdUWUftai2nT2X92RwxWa4zE5WyiIf3UHra8phH8BoIu
TFikgjaUcXYCgRKp4fA4bLdpeamy1Oj0Agi3MUAUYLv7MwZPO2+qDXPbakaz4p5n
lHDPylt6KilZTBBpRF0fZKVX1qcYk1LpmF8gTrTDo/R8EnF6LGJ29sgvVgVPsxwG
vTfrcXvZQ2m3oemPS4wk9Y4fdo4Yc3skPu/hL51JQPJuD+HWo8JzlCNF/gOi/DX4
TqNJDj6TZoj/68W1d8SqHfgUn6KCX6UE4tI22ZNMSdrC8pdcugrwc29smigME5BU
uLi5neiLzWHL2HcdMG8QEaDGiX5BWV1XLsiv0ht3bqgri5jODNoL/WC67iszagoz
s5WRZqU5JTWWpMjuGPl5rBftjZD+DOWO+jAxhZuWqaVAAJkf5NDvJiKk33avyELk
k3GeLz8gLqCRInfOCuMAs7J23+nBTfJXeeLqKNAERFnPcmg+P3MwLF7jkgyCKfRA
3BMZDRzXOl1FtTQc1dL1MUkozzn6ZNM1M9JjIdGrKdH0a1EGPv6PAkToKSBQ79JN
M0VPQuRjuk6DAa1OcxwVQWBQsWJ6PYoXcOL+OFSHxYAUZskjIWUVYBtn9wsLa709
YW7uyrS2GZi6N0ZwbGA14veb8ICOV/Sh8cM6pnZ7iAuFlTmBbaKRFmvSPlKhN0SV
jmI9zhA+8ZLbMg6yXB8lwR0pg0vObTsUJZCVwek9fAG/CUcc/3PTt5mPi+PVfW+u
/lbKReysu2tSTgnXcxLmYdOoy2Dn54/JI8r0YbtX5/G0NE0gwWI3tIc4KOWDltfo
eS1peU9ifTeni+4lhjdUgc/4Go9Zlz+g/ADJmW5GGluFDWmtxtDJTDisdPpx3Keh
AFMXIS2PY7mlQCbBSDHdmffGHysyr4dy+LFmdLcRdN/AvF8Ift7IMoZjYrt0aEvl
cVbFkDStc1KV/Iuu92g6jyEhhWsbzc00fftcQ8iuZ0PT5+2H3uTuh8/DhpmQvvDO
1xfBIOGxn0WUMUf3i/RZ+Ws8vXqaeDFGRYDE2OcYJ8QqDG1qeE+H3BSuJqd5tIdv
Ffo47Z2ZxHxGesnVfViIMJFuYGbFfVbgR3YpBmZ29p+8wZi95UypynSuFEw17L9q
gPSAugQa5URMw54qqwBB/+FAEjTGWNLmPFKUZs5esE0tpEcNsfChgsSfgseFWYkr
Cd8S0r1WlxWD9mZq7zroHpNodw6dSTkmOZXiLHcN7+5imGR2Ft4a3g8BsvTXdBeV
hqj/INrRs+GJ053FBlP6LYcQ0WgungbPMSsYmWsoclko0P6nfWDTO5IuZIfLE2Fn
VteZLgdSWHXWVTRmvjRPm+nZeLFv9IuCh3mgBcIYtqxlYV87iv/bKOY7KAy722VN
WEu1x5vaZn3Q++ElfcWrx/V72SDKGmgmoqrO5NjlctbMyqS9XavywOARpVgEKZLk
WPaOm6x7Ln1blrkrtElOWDE2OLdn8W4usyuksjbk/vWOgseJF9Lg3A3XsTA9Is4b
OJCfCdtZWELRJtMwJFayp/B88l2FDiJjEqBQvEnANnimzFBxpA3O8Q5tX1B8G9fL
We/C6WxbZXGhviO9KFTWOAmqWO4G/o2AK3dUvxcCGroKpJZPMAhAX3sKy9qWtIwR
OuWihafwoFbbrK/PuDN5GjWihUJaKPmlAdKRsQM5R5QLRjtnZJYTXV6b3HO70+oa
z8mHAHQ+PmEUriIK4kPS7SWrr16ot95IxRFHpo/cSEHsHbtuFJD0Ro8u8/m9Y3WH
NTV183bYajZSZzr0yqtt4IyFF+FVBKltx6TTCv42k1cM9L3juEG+r7ZLV8brhL8R
oD1iHR7sm01a/3D3VlmhbiTudWVVpGUHmi1edAJ/OOupdLWksEfG/YqHspYMsXdl
csmTibePedEdUl4T+ElTk21sBA1F+oYwubMHb9guvH2Wj6AvgLcA/6PxHuoGHOFG
f4eYBQn0DGreYynrTUXdbNX0FIZLYJbg1lqF2iogLPCXGu5otkY5LVC9JdNBBbb7
l+fkNC5xkJGPabjd/NaHUPof/oklEJnL3+W0OA2PBWnrsIPDPEvri3hX6eAu97au
1h5p2L5Gy5hTCQNmpfEN4zeTR6e+kv3tKq3eoDdWLpJVo9WekKKM5LIGgNCDP5EI
U7nD8F0vqXBD1T1JlgJ4MM1JUzpSBzR1FGiUEKTlrqcG17senKPctEyUYP7BB7uJ
90VBzdmU1cXsAhzYdD3+qPTUHPWicvayMDOdKZXR7JfbmVcau8K0TbeuLgMSgeTt
RWqtJqg7ZolSftSSUmFQz9sJTiBPYNKgXGasH245IsbqvCsM7UEF16gUTrRU3niv
pQV/DYXcN6TGU3XLxl8x70VkXhxVb86Tgb+4H/apTN8CgUYko96cze8kf1zPuemv
uNTmmCKDENl/w+zrdW4H827Fj9H5N5+5hAwZTArbQHu1/h3JwNksBS/fdm4BX3Fr
cK+ZL4bMtw7SOKgK0zXQbm947tD42KOlx8Ldkc3BIo+qknzeR9e8DKkZ4hM9DFal
6jOdh7ZkwRUx3eH5FEIWPksmYLLPE8/9ljrm967mCGvwvEwmxAgrt5DnJ6uYHGO0
bFBdmJBmCfQFcGXRzjq27U5lage1OUN/E+UiPNjvpoUnRUWVFzqX6on9BqQnwc2h
1zK1rU/IoS/2LeFEHWLLcMimhL4j43zInxD3wqVOdUmra3y8tP1tuhmcXNSGhaha
nf3xCOU2bPBch36Sw9KvGZ2EoddpUJDZ6bFIzaZhc/IJxZ3KMNt1mH6TEs7h9cz8
ezIaHPdpzilknnHkm2CaF72bTs5c6NExzYdt3NiW8aDC1P8lGsltn+kfcVL8LoDD
XTW2QHDHvvoc5vpTJAoZyjkw4fOf5Mf0Ro8JaFz6pxcu2mx9Sa+nb0EvYK07dXN+
4mDgElsv10BhzdbaHu7dJA/U/1gEijRH8fDQv+BvSwWbHU+sjj/Z/Y5XtA6XsYf4
IVk/ttYMQLGMU4nwqZ6Vw5gQqNjbdmgcF6WIblNzdhIPnEdaX6sucX47Odh2uzuv
O9tl8UMMWXLezC3bvVICMD+g/QsBqYJNCsVL1ulDZX5CIvLjp9ME+Np62yz/OWf8
GgTQ7c/C/fZD6GO6CXWeezkI+SdEFlg013Gu2NAWKcVdNL0/TYbTjyHdjwq7d1UX
sbpBiumHp5/OtAl+5gXcoozdOEAdF3FW6yYSMnnC0/cIts55YwE63oS/+JXUVXP/
9VCek60BijKiwmTTDntcMw41l95puWkT2F7qrkIB2HILLmP7LlX/wFlYU+CUbOsb
VXA/1htWdQu+70DNYTODYMC4hOEsCPYt8xDXyrI9FTKSqCWlpqCuKD1qjKwZix1v
njXP3/dapLmAi6QoaZKAnFAumyajRfAbmtllUrMa31bT2ILajIUs6050eSUu1oMh
32GHGqiEeJRJIsicSPDv8kAWJoWBBR9X2mhaDQS7uKXvSs0jLloLqSaJRKBwcxru
ONY9t08XOidiUiiC9bf6IVWXAXStohvb95hv7icU2K1PIUb84Yekw5rLZZk2trVj
vO2/vxrLfap15Ukh/PGDe6PvLjKBOfD0YuaAjSLMe4eVNP0kNvEVjtPx9pOzKZ9x
zd8e3XC+zFHi9K1WGYSyTs9hQEBhzkSVI9q+aYPe8IzeoK9U9WIvmd/lgAnh5TFI
aDNffQz/1WlwgvLkzQz2YKkJFQXrSZeU7WLU396qjRyVh4HkdLoCjmQtNry80ALt
8knKt18+yZ+njwTQyhiM2RS1YEgIHRJeCDkZ7gCWO5JddBufLCwinFc6BpCPjbPV
g/PHjYGtj4cL8NP8Ag6qqAQO4RudXqfiSNKAG3036ZttZBpTp/AKcjewa10rvKmc
jhSBpYyRN6og3XfcxH9T/Dx0neBZMhll+o6fzUME7Ov6emObLF0suldM3PP1V0i3
F/b/bg3+1SZBmTjll42G6jLRjS7n0sLzx1FH47/cSOAZVQN72/4ke522eKxcT9ie
4QpRETmQCFQIbyULn3Mc3hLvqWSBl814dqPGmoJNvQxf4MYTT2sm8yMz2iPcUg74
nF0woiDZc5i6VR7DcqCN6wgZdL+i18HgEKjnXMN+n0SJ4pjjeXBHg9FBlLkMlNaD
ZX57KU+zVcCkIr4neUHo+JPw7WIPalr7PFh8wi8l9WTlejq5fHWLGKxSGUqbMwQd
9Ifrd70jIUUl7fLJoABm5Om5a1Jno7va2cdtz+NBRIhHKsBaEBeqzEIH64mPdW2x
wOANDlmQPtSuRoyuCFyixIhQHQCMmTUzqalb7xQlnOx+zRGk1DJ9twoAZr2L5acs
s/Btmd73brP0Bgy5bupcZiB9goA+Y6MxhYg49GZTptE2Cs4LESJ1qjZy6Hl2mcue
d/8yb9tRjCmJlsLmDUfXQDzTr6MyjX7UQKVCqZ7QBRN4rlJZTlcblnnXJ7G4WnVl
sSkCl4TkIzGe/EZCekyOwNMrwI5u3of0TRQXJXmQeu95gITjfQvvCcsVmzFGUTbW
dalWgeSPzpYL13W/Vvsh1Qer+kzisTE41PDiysD9IiZXewDdT9DGCq7Y6iy/SW8n
clKYhEn9/Ts1ixYiJqYKpvtNHovfmrit28XVfBn9UpOnTg6M8+U8TdZ5BPWX4Hu1
CL75LIbq3jloMQaU0/wG9H3Q1Jv+FUgIMystEOzz1ZTUYNlU+YWnUcQbzkQ6SO/A
ggbg/AvuFTjr7mm2UZLVWxbchJNLy+gQdml3xD2G0pLK76r2myRHG9G7b0s/g4Ib
zhPueIT/eocoL1ZGn3H1A1jfgQ1tulMAZX5Of4bXX9cGKz28N56ef5USoQCgqCzw
geUdWBagk2z1IFfARTLWjRrhkbNfoZFHiU3E6xHiObdVg7LOzwlNjMNpcp/7H+A1
7h3EZNsyrHvQ0WN0FHu1NCaxvRe4xL4HyttnXhjNGSvPWc0U390+6jrKn1jwvUxE
UmpgmSrGolu++s3giQr4hp1snZpbXdQORFYzVDMnXXb5VlGo6865Mkwy5bdtySaP
PK8gZLw8CRMJu9z2GgL4onczDCSx9iqTEd2ySCy69KYvbuc8JIsuw9hFhphVLjtk
o9xnmg5OSzv3j7M74m3jGZ9aYfwsCEq4Sn02eoM6jolQzTend50vTvgwS54KElOJ
mGhHfzN3C7WeYvR1TBavyuCJfCOyHzfri6in/yxeduqgeXFYmci5McXIYTdtq/RC
aHSTjvTnfOlDeXZq92NHLcypyfkdlAxTyLrd3POglwYFeaco8xprMotevYU7ots/
ghYvkFCSzt7H6y0X0OEmqPFdi3dRRjgMQQHyor3ZbeWDY29LXZY0QW+xfd/AI2G9
NpvGGRdrSm2f2Es34SWjCoUgesxsJjr78n4Kmf7l1n9UGSAmYhoOYvU20RNgOfRM
ZDHkR4Id8n0R4Z1ARyJubndQf/36Kv0HRYlJrZedYLVAqZ8dOLIpVRMhCvCdhVvl
+fMbgiIm1aYOdJIXSgt7UR7uMv5r4Un0zJ1zA3RClDvVSGmlVzYf+x4Tmb7HSjHf
Tcxr55SQpVR0goCtv8M7os8DsCoa68IAAl0QWC47a2B9ohYvLYZ7oO/reRuyN4i6
/kD9KmsHxGpEwyZ2Jxwn219nK0GlzoYUhIYQgnxnwWTxVuk1eXm88Cvp0layAOrl
b2hsHF60PQl4JJNE3K13aAHRdqzyLt7FO3GjmOtXRuj1VuwqIpiL3jCDavb33eDI
Wsj/tBSlGLxMnihlt72B21t7oy7EEuAHb9L5GA7R5TEJUwl5yybNN+paMobFd0kT
5USt1IuYUIc20SK41atFF+gsKFB5kCyAMxS0BeOvePrBrJLN1LIypUeT6JA7PEhY
8HYA7tA+FtSpmPuuqSFNL+Izfi/GX2IsCzoa+9OEdeT/Ym9xAquJamZApnHLeu9+
8iLk6rX8hlkJ12Bw3etVQdqBJfkLev/y+earWsfRDLXhB1Nb8LxkLPs7uWPVtPa8
RPyEItZx2F/YdLF2lNgzllVb1jwySQtm+JyZQ/LbTHnJe0Pihp2WO1LTPvqp+iVc
yaudDzjAdnnSriNg9x2AwFRasy+9+lD3hk79MC3rWz5B+d10wTJBNkArOMw//jhQ
bGMHPkC0/9DoEiGEwjbx4nOhpv8vS3Mntse15VxS9BiQlWdNffiHVjpOJlw43HCJ
f2G3R5j1FEaRCiNOoGv3ww9/BlwOTa0A/RkGva0q+blie8eJYOJoniedO16HNbcX
SLXalGFMDhx6+vyC2M6tzEWeavQ4Er/RFcDkTPzT1+pyy89YRuFabzTGhCA9+Io2
KUH87o+A4vjvh7tC5xsd/adI2jrr/cEf7nSdB+d9xZWd32ok2BNC7rmHisvdHWw8
q9g2pwnqtDhu4uh5OigqtKFov6A6ppCOQXYKUSmFGbVtR2145paLMZcU6UdDQJBT
YgWAqL2Y1zQ9gRI9G08PEQ+JVAXcoOTZ2sKzuek14PsvthJWZVrrQriRQHfIjai6
NF2yiu7zzizzbhCrOM09CiynZDu5eyfCNATRXQtOA7Ss3xzGx73eVPkdqqMyprbz
qyIxCCMSGU+l1WycWrrq79wZn2CY4ukYpu/r9s39Rm1evzkdngYaZsrLPs40HnP6
RmDARwKCSDI7/EuWM86pA9khNJzKn0WQH62PG2KPnH1JWzRQQe34MgScijcA55Ry
Dgs8xig615IcybmqUZRQvg96nt5JwfTI5Rhv08U2VBUANW9AIEJdH94Y/h3CEc0c
yx6Z7yf+JFr4SI/c4QWCX9T3/efe0AlMX+JddgOY5eY2c99lAU8sFmNsgsd8q/c1
W6R1ym82436k8dG29sdB41XbBi3/RKbp5W7IKMnBzHbU+D31BGV7d8DjNtNKn9kg
A8XbKuqCmI07Lyiuf8TlUyaSg0oTuv/3vekXB9w3AorjTHuabpGOTQr/xj1vYAxr
tpdMMKzBMKmCBlHfi1wazaeBNox51O5xoYrCRiJxug3DlzMt0gVBx+GoZgireGxA
BC7UoiNUHoqX60yTo32OjlDajzaBEozFLOyprVqTHpH+3/Emb+PhNmIeEB/KpzyC
C84hUPEmWGfvKMaOeIzWpq0/GP/hqQYO8GOSy10Biz02Q3J+L8LRs9wMPFPTyETF
fao+th21tKFYKYWgf2RWTLH6pIktJoosHndagAh796EtGiqQLwdOce2j0mc2di8C
e3q7MQcGCq0IAUUybakLTC9hXo1Eef35TDJDRHiHfQ5POs6UjNIlbx1gqUdmZHGT
h0NzeqtCixzqrNqqZnJ2fVSGCU7HlkcD4FemtShQTy6hTuHvDAuSO5GhyR0T4Led
PjrXGk3VynySjXj38KlVgfEZtYog9037tt8SzVQ7tE7wQ3TsK8dodcYjjNVtFjwL
fY7NJwIAjCnwNmP277ZiC7UhTZPx7AkqkuWYs/gMy6MWvdafqhURyJcR35zaEKt6
0o/SbcxN0sNPLjhth5pHjkdeFclc96B3eHx8ICoQG01aYKqtHG4PeLY4qVGOyVqR
5v1h7ZPojfhQRpQxqkVn5jwU7c1jgQj/pIhWeyDqnu3MvNfxBiX+ewF8G5eCQr/p
hbqPtml1T9P1l/IaTfLCP3GBwRe5ctFsDoO/aywUkHljyd4K3/88QprCIZz463lu
fypKIVqTQMa0hzFJumU32PUVyrmEUJsPhtIL3lS4PhttQRRaQI7bWYcMRZQxsGka
xJXR5TS7lxu8XMCBXuhCGtAOlnnqRlnR4GheWc4ItbNW4c1jRzuPhvPPrYbMb1zD
8Fqoa/WcO2d0HDWS9jHzxdkqXHSCJJ+pJke2kXxpKkesE/0017OLioBWM6fsKn/s
DbxyujUQDdqzXoXcZ+ewiaYJGxgr2eVJdBlBcqN0rQU0BZWvI9PVlwgTsgJT6AgS
vsNnAwBuWpbAyfG82VqttaaOEH8RMBYuBpnDOb1eIsiYroN1qAhmR9RbGCHQPYin
RlPtzXHKCspzXNI1mtHEl5CWUMpZfSftmOyQRcGEtHxEmIte5Fjdv0j12QqCBnBY
gN0wC+ivhbYuFErwhggisLjs+I2fGp1zwpvVrHgge04Ycr59nhisV60ukhsJbbUD
WLCOtnwiDPWo52oHODjOpIQ4DNEVmyZnc4UqE9hFWv9AVZk13/+fgSIDNcG71zmB
+DDsIRWOklN34FtWbi7kchqs0vHGTtBMqVOIWRnEbMao23omQM1zxha6YbJ1REyS
2Nj3pHSyyKhdctDCN8nxvUWbXIBK0+sdgUd0fSrHbDwFuLhpI4bUF043S0yTg2fJ
WEEzzUQvI2tBF8BjZnnSCtiNrdbjQVooTuiB+TvCa8pd4JAzWvBi82VaZFLjYQz1
grXeuVz63PiujoppgN44JX1/cPaGT+xAnpyv8XX7xkk7O+J0Vo2rZdo9+sMRdBGR
l3H2355IlQEdAURMP0f5SCnKex9+/kr0UgVKr+CQePIBDK+tYh6KKlXaHASPGRo3
poETOtXU6+8+PWWZPvJglil66KlpmfLz8w6j41C5LS+0UW6pepRQX/1GXvVM/oMc
IOSBR2s82HwRD+l9Q8xZUcnBoLvQGSmXMce+aVjR8xAw2/pWqFbF0PURxk0tZdsv
faqPlLGj2nCFHs7kVJcN4cW/bV9rKCPPWxpNd6lOgfCQ828z6cyT1V065/1MkIbx
Ufq7WFx4Q70K/mA2l9wCNUPyta7imAEJid2Q9fl8Ied1j2ACx2oR6QhgQ2pLJVJf
YdCtTv462mEM7uhHzsBVv/lTsc19HmdK1movMjVPApFiZrhktGQBgk8mETEhP/My
2iQ5b3G1iNoUDSBOJne4orGKmxmTd0TtMC/6TRRHpBEGa2nNDjF0N8uLeXL2vhqO
KFyV/hXyh18M76HjzBikJm/aSWrALLb82Db8/eWjeTNHjk1lK8s2K+4FiPDwFkNu
xa8ZUpYg1sh1Ad8K29JOiCQg69JDjvn5ZqG8mlIsZLSbqgchY0DTZE2ioMZnTpbV
R6PoAzrWKN8/i8QUfFwN8n6M2Va+B6hn55XsDUI6tC4e+fFWQ+9uoFEy8ZKw2hFA
4gWck26MZYUWPKg7T/ebv/igsnQkZV1y446sibSNWezAkOBl7YdyMnUUKL56L8kz
x2QHEQWBhJ8OpHw1dlmh3kFZndHUrveluhLz/woVIoGOrZ6r0rBnUfJqmdI1P4Gu
5xUvGTpn7eaHZjiLMtxdFEpNAEAVz8tlNlIGXw27Quhbxy2QR0kOLZD4NRpHlfMk
QWJN2u3ljvUYhkWRCHhX0EOrvKpkP63CwyCB9llRh1T7SFezaLUrU5laDO5wuYE1
0XTfHUY3kfR4LY2KCjN7XyIOtVEk7WHk9/8chAgtny8AFfQomq9eiCsBBJx+nmaG
5kM3Km+Dh1I6f8btMVi8CH6coPZ2tky2RwFP909uDmeEMOpSq/Gtgz0uSAAsfgKx
vNVLSO8Z16w8ZPlGcsxd6VGZIbUvc343HD86QDt3lMeZgK2AZuWixVPmHT8FSDkG
huBZEHk8qhtdb3lHfD9rNROwo4BgpystQ0Yd1lAts2ZNKlTlz/rkyIOq8MjYBl3n
lE+JllzKp673o2pIBsA6hxF4iZNDdOdRvtrCrx4tNkhewhVt4+k2grXhwwlrRu90
3GKa6Vzd+yKTgBtdyvYzS9LB6VESgKh0Q+XtdPcnwsPFbJGwARyFE3zthhns4cB5
6eSriV85XROzc+AYAIVjTCsE/nvXflcGWEnHtKZXEe7SIt4JU+5/62QrTUdEyOPP
CksZktkK8dfNqD1/nu/VtaFvoRCyY85C8Ry/KwCxjdtkmIfRS3C7vTOE8KLPylxm
o79kFT5QcZKbqXuUHe5PzjvvVRAwjT9y3+9vUPfpn5d0PXJIKQuK5Iuj+Am/eZLK
ccd0otsKGezCR2WKtFgMKezUmgwenxuuQno1Bi++9jafX47HRMYbf8BPqCFueVqL
qLSAXc6tlzg1n0CCleNhfqKKlezdYZCzPdxToZXFzDeYBLyjkcB9o0KoSe6SUgMi
Bam0Zu0/k6njd4aBaqkYA3OrT1BPqUfla3fX3d9CSplOBw/hhB9x4C1Tru3q4jua
tlSao48/VKd0mHaCp296BrLQM69mz50KMR612HYVGMfd+RvDsnDFIt12Z6OBsj9X
3a/tlQTFKoLQ2RmRVxDvZi4+YuXQwlgFNR9taMyP2xHyjuUfL1IxEyEItpSuBUKq
us4y585nhBX98DUsrGI1lmw+neLlHMpCDDAa7LrnD+5xuXP3+3cRyCoPParQpFsN
JrR4yle2WSH40QRlDd9c8lHpavo5gH9PblXtkdbolL3+JtweHAu+c+K7YOpeZw91
P07hgsV8Uzq5fHX0vu8iiFlole10spH31oNWR+s3evKGHHCxa/H2JjNe6NixuxNM
wwovTCEkSsMfXbvsfysJ/CX2mWICQC5kiZUtDVPCcSlDQHpO0VM+KjHjfyoMrOSJ
ipI6FUiREYxGC1CyGSqRNxeBcGjyI2zr3vnQpRVhQux0MFSexH0xLgFbrus/7arn
3DdQycrJuWGF/mpyi04eeeALqaXvlp6wLKfbsr4HHYpoG65uwZ+j1A7sSlAVrI4i
IOAdvpcnbMHTZFUwHPIlMvBUxAVjKJiaU/0dJlTl0uMJpOah+8st7864rFz8al00
qOB0eZpVK8wZuDABoyb5S5S7TCBQ1ECBPFMAQgRj8zV6IqEJkzWGTCAwbh17ZEIT
3iXUgih6avjiqi4nStUmgztAh1KJWLiCV7QntFXbTJ7UhmujJk/AJwYKZRBzC+cP
Rwtys9VWlbVfQLbOxInmAPEx18mNEdV3p9JLsLD7zqLhaqpkENcznpgKUbl0R16F
68w5pY8LFxxclBMh7SKXvv2SwA4rMTLaYpZWJ52RJye8BGzzjyOa4h4zcvT735pD
+sEBegCrXH0jkdtLjtzRyM6cj3CTjPAHMZYnJ5mz/uv+hQVk1ggXlEFKuKaHYdzC
hKMULiLSMFWj0kKqmXJ6GGU0Vmd5rSlaEoplEJt8n3abKAnBCrhGZLfVjE3/Jk1a
g0X/YZ2aA4PPMWIC1tOZQvJ887b4TLMmNqJhORicp9xzuFnvyRJ650gd2QrE1IaT
rxQTR5CgsCmpULTTjCIJ0sUzUth6/blbDcdpfmKQke3SLqVGFiq6hmNxssA9DxeJ
aoVSGle5Vv+JIRrkN/pZsRkaEa/otfddXWWz2//CxG7pzVQExjEd7fw+Fse/q8Yd
ZgUcIugH2pe8x8A8Cg4VSn+LhuCBny67Rd8a7BJARQ7mvhh4LXP7WUI8+YeHwnLY
R/VtSg3AUrFMFmfUr+xhgGadgMMrcMU/0huftMUATBkWWpX5EMcRFENP8fer0Za1
Rftu46ClC0bmg/ZScHRm0fz4xAIXgVqOEEop8Zw9OH8PjMPumG23LlLPuRhVFHb1
nta7KlmXHej5mnGxm1o2cf1p45tPH4VEJjTmqZp8B1gXmwH+qPq18VfgC+pqarVc
adJKPFa6RGx7RIAZsTYdYmn4XmXYzC5CC2Q+6XwEXa2JKMfTeIWyaFPl97CzqrPF
ihomC/xYQX/Ee3v5lMxBQkhliXS6BPd5K2KPqhPIPkEP17bb12FpwAu4vn9kMMpD
w4GaERqvwRkGe9xzhud6K8h41LNZXPOU3I6+iFwZYciagAQmkIoy48UVZ9ilYyIl
d7dWIDwDdu6RTP0G6483foLHE7xNKtRmiWqbC/XsF4Wr7qcuqdwliidOtBGrLGA8
ApPVjiGVYlF4wJrx+aqOTVN9wzQmTN1BPOFEZvHpUy9cQS25dSl9YkHt+ZtXnRRL
YW++wBu3zH7pfoedK2zWbuzAu2Syx5ZWbQAlKN748EVtdni/1UUGKkWu+KNVPR6P
9XsVhLMCsmtOi25cDLxccPbQ6cb+hWGDQpl9LM5K7Y8UecuHtE2PpEDSMP91oA0s
lMq+VGE7A0fkPzGhMQ+YNZ9SbCSg/BfOIdW1JZH4Y2vv2QrT/y1PGPPy8IDaXniO
mkNtCWCYvF/oM9Bj0s34SR4oDwTgyMvVJgQ2u44A5E3qlSUHo01Ft4Q5bQtArIdV
AZbBdu9RctR5jE2qFg1/MJ9iUz60Hlm/Hn5IhpiqWcumvLQW6BDEV1e/PbNFfQP8
8OfO4macqLWjkKzrqdtLPTYOunlRu27/VNig/dzRP4+a/fNFeKvRp2PZcK1ZjF1E
1x7BXaOB4cPEsS/X06+F2KHRpeOhifSoJOpmcHKFqOSZc43ZzOq5h8g4SOX5/BUP
CLaRChakJXXJnEyc1PoxngGCsFGgQJvrbF+MGXp8CfrPGMKVy0S3qYNlTIznR8hj
9byHvC0WXWdbjW8+iBq69POUygubAbsd47Wj3KuRXO9hW46Uv5Wg1MFCCxXHOHZu
4Ry2V/TbVQGsfrPwavKAiTnaXteuRkz4RAchWCn5NHKAvTMJm3HnkTlamlnYYUQn
4OZOAxuBWMFLO5OKLRC2NvDvCmW+bbuS6ApeUWQiHIM2a2QSSa4s/IZc3NJQJDqU
GrxVm2JtHSo9AoLxwk5ML13E2Audg5/wvh0MAKKCD4npTXWwE0eoXvDl8CHTum9B
5XTC71/Wy0QePWW2oWXk7m10o+n7yTi62oxS4Vd5f7sMXJ/mgc9BUuNA21Lf1q4/
pRGFPQL+4Js6bKqEAkjoPY+lJmfsVa3iWyfbWloCMV2EAHRfz1j7Or3AUH2+PFLE
VRWQt6+z/C9hrY6+j3ac/FKZj4NP2HVoN+ny9DWh9jiAvvpp97h8DdLxPeZI3iNU
RjcQZZu3bJG0VgHIRfR2F0s1dIcdrpBQ/PzdoTTFuGvpJWndjwpa6uxcXo2t/NM1
Q24ItvjNiGn8y1wVwqdDFCzt5hLN1I4k8eOFGoU27KKzei9Z5E4KyTZ9onPJxy7U
zJDl+gKMkB3im7kYirPnbNLIv1+RNn+cMNYh6v84mfvnSVDF649MWGetrM7B4hsn
ZHNAoYcTXCMc5M8Av2lK5aFObwRw91G8jsbDC+6XDIgWDswzzMtJTnO69SMH0u3G
BbQkiyHjYvMOOAy0cjUt5D8DmgJ3p46SIYWdv2m5WkE6mJHVkClMASPOT0K81u8y
f7I3HlwnQ7upAbTbn3kIwMuU5DuHS8I3szJ+/SpHtiS23FQVY02N5tlxl0BXc650
TkaW1vcqJicgxbsZXKDVKCqiHsetKlQn3hT/OduTJ7oxYUoP7Oq2+4M49UgAPJ1B
wicBMshyDH3a0MUAdDgyFgHJB03PnWCktHD+t04zVIOR6LllPr+g9/BpXF0HrzCI
5gADvK/Gw6Sx+K4wN7MuVPQSOllV5HhPPZ1Dxlh83enmAavHDotTRsKqj5x8nL/0
ahAvey56sLy//PAS0eEmgEZGOcs7trtKZt2MqvpQAabJPtEtTv2qBQ9dnQXbThN5
OSefVpmaf9J7MyB6VGLPui9zpOx/OW9ONUcJw0ObPX2Y5+fm4JDSKRcPMl1Vl4dW
hZMvRZDHoot6ZV4UzSBVOJPIr8fx9kwxDJl1OjKEH4zgMZkK/geX2kMPQVUC+P3F
+aixL2bMLr+iDAVphmaAznK13bblczzs3PQ2rC9tmKcXg5v6rz7KMvZKKB7TUwhC
P1BM9/hmyQXOx0sPMoDWm43wlXc4wJswxJitDk1BEyQl5JPbvyhAR3Zl8f2+Bw8u
2ZHk4DaY+sSAlocecNpi8gX/D2mgx0herdlhXE0p0aj2qddPv1jeubLlxKQVSZyt
UwZI8gqdKbvYYkTd2eeU2Hr5qwG8eW7QwVoHRpOOc+sYLlB8VnrnyKP8BlWpsS49
jk6AZHw/omsEkkkudLu7OifzALw+zEwNhw1aKhtWH6lydfcQQX10I4BeBEqxoTDP
/UP9hcS5O3Psolbm8+oRLPgMOJH74nb7fcWxYcnSkMAb4IahizGBGaOWwZ3xIjwq
uaFEdN+b0opxy6JWqAWavtXRZt0APrf2LdyP26q/+TmNYAeMfyv3PPtdX9o/CU3S
YGHWCgMM+GH/hgjw0lQU4Qm4wqe6yj1ciMngU9ZWffkeZxQjx/HBppx2uycI9E+w
dfzaO1wEf5mveKnoGhfeSu0Y8KsdALWAuNVe/QjwRUO3rNQFJZ+DmZ6TVkhlOqyx
jdSYqTA5jAvLk8+nA6YyUhNuY78tpEGEE1BF7mCmHA+kwfqVHUIxirD9hZ5A4C4V
T2t7BByVAKauwrvRx2qt4l7PRkDjewRADb54Rq083c0gTFnO3JMkOmX0JSaUjK9C
aJPWwqzisoq4HPpDwfsfoOsjDdEOx4AyOtUqK4zOpcQN9O9vg4J656vw8YlxamO8
+oCz287aVQz/gorYJwH0nDfLy7TqbzCzJjgvSaE/Po6ZmNw1HdJehkW+pYIzCmsd
Ra/U8Js0seHpLujnowcjvQ0FZ6RKbhauF2yPByAQeQTMhqyUa4KxzFTTs7g1/89E
mct23sv7mlpLUiajr+JX7FpZohyIdVb2aBNzGV1AdG5D2SOaLLvaFJVU73yM9IxY
71kIyWjKRUFlvSLmHsxbr4xJdTVJkNnH8sLMJCpjZEDx+zYAGFlV9tVMAhp5q28r
VWne2dwTIJezj14t4/JPMBjVR64wuIzNI0XHEHEYA1Vzxvo4+UWfkSU8BR8ELU6i
LkbmKziRaj+iyt6+Y/+Jx7Xpm2saeQeYlSEoL/p6YFpa3DafDvLQztw7GIwj5PgQ
YbsRBHiSo4OESvZJ8g2ggb/DFu68ZbNgK4wv7arSjwaA5nS1feLkKjkHUaqBoeHH
8bU+7YQwFOShLSqtvKZUbP8TCOxrB05pnlIndtK9jb3g7iqV5ZUZkexDjoP0IU0M
v822kG96Z/A2t+DROzknmrRzKM/K8U2i9u5xJQqCbRsXftLkvZl776C8KHU6SQvQ
OktVR/y4ERgGdy6+mzDB/jSMAz8rvC0Gczx157ct7DjYf0HMnVoo6zUPdcIjoT07
SeKu6GVbavOefFBV81/UL8CidOJ7YhvjOwzHa8QVoyfXFvVW6cLZuSHwefme6ckn
ZDgzGjUibLiz2OEofmM6csCuEV2jaG0sgiVFb2Acf7xyKj2wh2E9YkrLJy6cj3fj
Op6eNzOERhj6xz+jOkMKGYQNQUK8SWfxr4m1vJDGiSTjDHD7DP9rQyq7ZQe+WYtp
HOlwuQKyv/QLxJuqm7cd6S/sT31sp/Aoi/jZqoeLgnUJzNszDKXZ3IiJQS1YZv0J
S7ohEVbL88gXuy4OPrkFZz2DlgJ1mcBmsEBZGGjGLFQK7VHb4HbH3cFB5ftAdCs7
w9anR/FNMmVJhroAfn0BblUiLixEviBnk7jomffXF0kadYt2GJyipTCZ9/cXrwOB
2wSXMR8wBfK8W1ypPYQuOwDuK5iyfRQFZQeik1S5oiIlYiq8ofL5JzRDadvzRw0O
7HSaIkhU1BwNQpO9WUt+cnr25lM2ojzVzVlOn8HPPgOdWGO9W0VG7TIGK+zmr5sB
MdsdMOi8VwSwDRsn9cLZVGAaaE1bv66xXJGCr5RVlIgRHpsOr7xq8csHYlgZ0q0M
TAI338e6+wI4W2sHTNfkkiwU6tupWDkZHPePnwFDjsEjmUJMHTlgoPkoFROFPRpC
Oo5YMMLFBu285r9ZkftEZY4Z86iuMdhsQdCHjeiyALPy5fqdrV/D+F/+YEczpO1t
jYJLSw2AIfWE6K2rS73uXi8poje95VLZqOeHWwSLfFwZ6eCmH9oQ52/h7DJOCbc4
bO2b+9jjwSR2pgK5ImwG90JoPIWrJUZ9tk3eDvive87REnu3FBVpiLgm0dT4U/5U
htNQY9aR9pObc1+T+0jS8V8SQ7IuYVWADSnKvsAkPowOqpb54JN+utQtvXtATqTK
Lhf5FYSxfWuRU5qk8eowe26FVK+y7/hKF4/MvqptenkXWMDP9/Wabtv801pxCQ7e
dE4nqTP9IGx3e2GhJ6qLdFYsJ0zReEsbWa13hPoXsTz/IuKFhIjmAtURgq8xyF4H
BfHa+n7DdLOPSHdceC93umJ/hGz+VmeFny48tsCHbumNm9sL9JodsVRg+VtK9mQI
btkmDueu/aFZJv+8tectse29rDDs45uioCKTIqEzJDWWIczlX4d9bFtbuL/StRzX
pMcum9TqAL6x+0ioXRKYSRRMhUMec4kdHInCJjub31Z1ifp5mjTaCFf0iPIOlMpJ
4gmw7STpV1smuDZ0JBEez/xyj5O6B5LMUdeSFr3uYZUEkSn1KxCGwfRbKDc7Wvjr
PQHU4f5Pl30tqZFzWe11E2BPjTu663808APnJItlSeUjh/oLZcy9TwMA59c73EFd
K10yF0JZg6jt3jOlsCdyqTX0uBGy3Zv+x2SVJLTL6VoelxcytSrVGIRqsYXK7HpH
mZvPZDJHjshKTtZ/vUXcUor/QlZAZbBIHoFvBDMO19haLYqy3CB/STxav5iA9vi/
mlK0iuJ0GSeXjtC7MvgTzdyvymz/G2RyFj7nHV22X/TdVU8GoeVF4DnhI6cWHPtU
CME+gHuZRdlvB7DsZqCo28uDNEQjr3OxxZlFUPS2NFraVDtyUvUpGDERwfSal8JD
RbOtGAJuI8ZUCC1lpamxsSxYClpsMBmNHyhbAlHAmatqv6tmSKVApr6f2Xv8KQh7
rS3gjtgjQVTR1id7S82dpPVOtVuTil71O0gSFHInN3+zMXxyky5nxFOiDANUphpO
QbzEkMAJP5CmV0gl+WA80zxkQazgpCFEDW1Gy7XdjsrmYQxSO0bii65HISlB9mwk
11cEvrKp0pOUyzo/p+Vr6SQJRD1UpE7152mkllKTMw4DhpQmApeT513ioXquB/Cq
NN5X7oCk2DpmKZABCWhtww1G2aCWxL2t76kSqf59rFmu4VOyN7pWpN04hVcg88yE
fgK5PCaQ1Np7zAezABlqm4oWeHK30fIn6v9aUezWOpGdHvUh25lrbcZK9FlqbjXI
YdlK8y7EhHwz9vPE9xYBhczTV27KsdacOpAS28JeuRwscaOeZR9qb6gwQkxWg9ti
nFHBw3OmPIVpnqfgQCAMDpCtN0e08hLy8sUhVZp5Jq96DHwsTtlruUU1zJd1WwO3
5preC3I+EXhM83rWs5SnhAADK49nahc2AMht2SSuw+Pn9u0zrIr249NRIDuN7XBv
5hRE6VsZxT10WEaV9t7SWUtowRQ2lZsweW/+bOCq0+DrO71+gflTJ1iT8QcZodKc
l7YckNLYnGuq6kb0rTMTiPedM39D4uncPzVzf+zMEsMYzsCPQy0Y/D7u8SF2POTJ
1CD6sy66XPbiNSGhN/7LyCPKNeSDWxQ4GYOPOFm8xa/Q4XxcjPCvJJ1ojHE31MV/
lSeWMIykSVvzIVU8/A8seFPpop6RET90MfaW0w+GwGNYqhBa4bYyr4V6ncdzv+/v
DUYi7eNKwDTYJlLhYV7otucriK9LPr3RekdJdCiPm1YJXmGbPBjWEBuZCRvKJ8WZ
04nMEIb3gxTLB9rwfe9c6uFzp5omks/BwQsmIC1CSayAazLwKQLOMcq1oIstztBx
XFvhE3tEvJsrRHSvVPZCr1tnUZ8/xsV9taE2RyDd1UeQp3BNzxmAW2qj8Xbq1zg9
idih24ZnylTLacOILovT7qcXH5ZNeANsJbxEedogWwhdZrPFgHwF617ClnmA69A0
wtV9ueYZHRwVlNDwAHMkIniZjMT7RwzRn2Y1VojtTKKy/t898a4D23MaIm0+G28L
6qYWKAbR/IKIArm87VEdAC2Pt1rmXcj+3WM4ofiyY9lMYchA6ReVsvW0Cj+07VwY
pnspzNXJ76nvuDtvBQCFdmEytOZnQxYZHjGvY9V+UmtHmhtZtJT3l7++6hW+sfRt
kl4+O97dzJAXsoTB82bnlIvqnUQnxM/15O1debGEoTpZ407sJ+IEg/3umE46B+Px
rZV9RsRCKpFZlDvJXbVnJV4Nq8ZLH8Fb84GqsMIyiMw3EpKPd5CD2uabEkUvscq9
up07E9xxZ0ysDfiO+zOuy2uqPDri2jsBApAz2jN0u06y5cxKdvpFurrOqaO+Yu+f
QkT5YC2eYTFHNqXe1vwgFgawuN1tg/FsujfqYGcRU1NJyIzDp/RqtxqpmU0NBek9
o/jsmSwxZoapgfWJKhWyI9GmoABQeHbnPR6tVZkUdB/eng80jnMQxCSTNlm8hNuD
Tp0BpNPcXOAXHT5vvF9MWjvNWo5A75aMsMajYr3YBrBFb+CuevRq8Ni3ICG//sTn
/OXvLzi7Dw6IbdBzY8rFKDASyXYgLW1kjoopXsS9chxkltDwzyJ6LLZBGq9Sktaw
sChHCT7frYZOgibdig8+8mONMvhoEgwpHh2opI0z2CWtBpNI1QJYXAW+b38IAFGS
xx0ffEwbL6EcdLN5BC792aJo9tf1UTd90XjejEbwbshwVIUxRsPCOnrrrBjaAwS/
jOpxmtvw/457Kq1FoDahVcaY6LFR5SrHT0p7t7a8Ekj1kTck0PnOqaR6ZJsSn+CY
bnBpyn2AxUxDPy/wbCzqcInx6OB1CGRNF5sDJW3bAUwG/jNR/M52wSdgGSRrcwFa
t9fyoaeQI4a65n1HzO3g/wdGQHtRxpva1VrWhcdj/hVdiX34ukunX8dLket2jvd+
ASLDbF17F5ey7792ijYSdEXh789R0/I4G0TIht5vNVf2PH6PBDxAw224wV/Xp5QJ
BmcMmTzHPqVvr+889NoZD7t6LRWTqDWCMxKZ3TxFLBY4M5TDWNcFlWiPYbWI3sRr
m5ocXiRy5LBCdiFl1izs5hbAwqBi2BYeRSs4MkFJ1/ohWAHSLiNOE96Tg+0aFDhi
zhmoaxF3EASxBOqPkNLnFWrkUoCd4TGHYiJai6UPscb2k6RlW3Ydt/oAdSgK7FS+
O/uRfhmbpR2nQo97qodWobHXJSbA/7fc2sx7K5nU5Ed+NJUnGWqwL9ZmIVruGQBx
d/Lzz2b5/ae0sb61jEGSvJO1ry0Sy7ctaWnTtQngbvCpLyCrXrZkiFfguKjUJ3QX
DSy3Z7y1m9GuIA60uMcz2QypsBpz8cuEdeo2ILv0C3uQs0G5C9M6CGedl+0sC1bR
ND4/zHJwF78fdKtjhIcaMgLUdObBY3QKfzzT9g7/be6sEJe9oqF1TsR8ImNAsvVe
K+fTvuwJjZq22AUO0qg3kFeFCJ9tKtZiMXz2xy5N+zaWa4+m0qCO4dKLmlWdxFs0
ap9bZdCgSBHbF4kdWHPVClr+WbS1kGOoCR+br/9WhhICEyVw01QvuMBscwCGh1CL
xM90bdcw0m4tBqLKYu8SXbEchqVPtUafyrT67Uh5C+TWldRFk4C91StMgO5Vx6NG
/OTetGDp1VlK+iSS7RxnVcFz3vpqRXemlN6Ne7HzEyP0QGkjOP019SMNUzmdwlSZ
e/+Ti2I3dUDUq5dMtBRs1d2S6uPnszzCS5IFZpTv+fDzNbLvwx5T9wIk9B8GTRWy
GSfQxID9Uj7FL8rNUr9fNH/PGH2nUJYOAWV5rJJZb1bCEE8uMgSWFFEkhIVfoX+8
0gD22WbllsZSnXbvoUMrcN0x6NAzv088s2p1tBn54E68nkwgMu3UXbIEvauBMh0b
D3lTHokitttfXzSySJGfW//aYuBlpbJ9atnX4VZGwiTyzHUeQRzyvpehGdU6H0wq
g5LvGwRNVuD9R25n4e5y1ydK+H9QJ7RMH2cItLpEGmp8Qkgom6PDrVu3XdFAJEk+
wvPGgKHhLmgjEY8HHrrqnXaCip7zRwgVJ7LJoVSmuudXHk8of7sm8fv/UqxFYk+2
AtcJQZzVTYN4SdLZJVahqwv542C9KdREk7B0VC6shRzKuXqqAMk/XjIvGQg579s8
Yd6qInt8CQ7GCRNMM2AK0beyVVtRniQZdmcjYTMWPPkrq27TZhKnh4P2nywa1CD3
lpKJ8cs3TGcU4Lo+oWT10c5C+ocgHBi+3yb4qRdY7O5xY7MGTzFwHXXsfN9bDa9G
9tAbp1BWW/RTOQQIjjCmgqwhRB/t3v/0tCJldJDlv6pYOAYHFRWbICvgPMAiGCEV
pJQXZdhvZQqZJsj5RSIfHzaGqK9J52hFKZILhNdPQ6wzG7VsVdm97du0CbMTRtjA
29ZV/MJmAPRitW2si2yVRQWceot5S5xidVASsBbaAOdBTT3SShZ+vUKOTt+qwAL5
DT/AjFJOezZDEaFj8Y7Ix3K3trv15oD/KjAkPiA7avV7iu2QOjdeGgQ5WxIcXz7Z
RVEnvBlLRtF/krEUPY1lJkwY1sdXrKBR/e3l6fDpx4iuuJbiV6FTpFXErG2Nh7wb
No01apBxR14aQUYJdzNvoiDdGNsHfypYGxsJ9lz2UvWIUW9AC0duPIghzaZIHQLJ
2xRs+hJj2LEIJskqUpQo/X/b3YjEcsmiuKRH9fvCWyAKuWHqYh/FkqKLR0bIlBxX
3nv0IAkyjlGTDdW+dxW8LySftlwk30Yx1A13eQG0OKZH10r0EBscEEA/atBBq9/V
FC+rRLr+CKi6uR0R9ACPYlqWcAuEBoVVlP3qbgPeTmR1mcPCCL6cbBg1qYrCapO7
kVIMhECwS87hg3lCc4d4O7MLT+bno5h0Kz7w+7xL0RCF/5YyxRH64h38ylVXQ8cw
uEV4X9wg98ObReAXW6vN7xV6dmYGRNlFkUwUBOifti1ZHH59lPwxkzqLMMaEFny5
965zhNN0aex5JF57jZ5hxrO0RIlaHlsM8V2x+IJX9zUqKrEeoG6xJ4pjjg3Bf4IA
caibJ4uoZ21HpG8QqzEOovx02S1sTx2CrYeBXmevmOPZ0Aan2BqLjbvMtTfPdJDg
U7GeWu0M6X9TCBgf8/pARfNH2jm9BNTLd1H8vMEDBTAjPF35Cxpgu1RbyW/oUP80
FwODkTFjJkxyZtVs0T/91EQiu1TgoAQH5+y2UAy1rBv46NCULKgAOpsJFBTdNlkL
Y1LuZ5lFb+baTEvdpjWMWpxef6VftyBjYcTkTvpTpiNrOn4491R+KqTKf2uKRiAY
dOp8MU0hF1bcf06U7YHCnAMDMsKX2Oe5F1CNDCpIGnn5I6P5ZguMYW4tiYeU4H2i
BpwytTg8Kc7pXqBEGAjngjz2O7k19kSHn0mxK6kaOXqkqz8IBwqUWEkAqPh5sBS7
fxtSu4toWUa2k0xptGHOCtipBaGoVJP3sY8uDiGppjnnXx2xbksF+vz2eR5vJfBe
IZ3kA0UHHGc3JAbEoCwP4yMhpSua+tM4wFiJBkiIKZNmwYXwzFj0GKHIWs4iFLgZ
waqn25/id24mc8N0INh6N1NUt4I5jO2vyF79jqPVRHb5u37vlEmdaonwDRHiESMJ
xBTvigEYBZe60rCoqP9cu10Um+9C/XwzfvaAB5Xpj32qKqlUygyP8tya2druVCkc
zU0a4nUau9TpaBI1aHtBJIaOnQ6/Z4tidh5OoPuit0MBHTpGw4mgNabG+riUtlef
BXrJ1rLJesm1+cL4N9eeTPjnLpxFGmqETnOCk6xB3ol38KQVdg2n4yBBCU5pbHoC
OGZq6zMVKLtoGQJhaExf6XYljnvuAAjcXRxaU0s4XrGQixN1B26b2ts8kBbpaMIV
GhBHjMZcE4j1qI+VCy5Zsk2qHikuHLNTL2ShID5FYG3ASfmdlxBPhUt9Qe9CwWHh
k0tTYhyQhoOWj/WXu5rFqPumoc5dwzoGMvpP4I286oPmHwka3d6bd5IdjEED1r7E
cw9oNjBJH7i92AgsgB7i+nAzlcJKndckMCFW8P0XJF4lY1ftxbYxrUVSK4wAFzWo
uLW305WFTKScMWQ1D456dKUiVOdA3n7rwGvHmW8sBqwq82LUailNV34Hb6E9AN3h
c5SkPPq7oTLljcMmYyUgwGnDkXtbhJ8RD9OjQYkWuduz6yRDkGCaTpG+MoAGfr3W
y6l70rZf+hb9JqCx7bsBAnlNFTRkXrnpVW5umhMq46s5u47PkLEi/5pzF7amBtoL
WAodR2FohaJblFkOMKvsb2yESMIGAiK76R5wmizI5dgPv6sFBx252fDpicEq1twC
iHuUsIGnpycgaHWGmP0uOBPDjSij16u0vY79BDSL8DMtGbtOdbWiXlVCos2pYRU+
TbL4YNH+6FgkTw5T0hH5P7M02zcQ/v+Ma6lFduXuYmhgPKzyKG2PqXtymhRbz22x
2IMpDrsRfUXVFEvLOU3pRNTw4wlNglD6bDWKqmrco7owte2auXxR416MWxPF3XbN
dH6EDcIyHlUHuutQX6mzrF4wAke98hHwiJeRBgNOLi3Zy0p/oztfaNL4hfrr2QDq
PjjsqwhLr5gdC5svfFtGnmP2UmcDod4SIJSqYv7DUlJOV/4cImIRqo9PLs3C0M4s
G14JZtrGfwdoDoVo7LiFUvVHQBCvT7GXQuoGVDwUxOcBuin4oAQOQW8/c/ACvcCf
pRO7NEUIg7fRdc9dANiRxIum4gOIQsAnU3o2j5jYvHr+fj05YIsKJuZaJX8HTDGK
SFTtNaK52f+CZ7AZlFRlZpKT5y/XGuxdEKryx1Uuac5x86ZqS6c8FY6cN3DtcW2a
W7BJtDUfJitOA64U9WT8mI6qBg5/oCj12JEKG0HJL9p2KdAVtSemmp4aWuR7bJ1e
4RtTUhsROXtBiKEn8Kaz8CyPQszDF/hXv5B3hk/AqnET1nJIsYYPeXJC8G7dktjZ
z8aZ7rGlXioFTy7LxMH4ssXkzvBwbPqWDoZdhphAc6qu1Eo0RQroUDsdGN/INtDA
F5CNKhwXnW0biyO6S/L+CE+D714f0naphcJrL2XjtU4hnx6u30ijQr3z7KooaQMU
gi+taAou/223YUNJP0X28WIwSM+MzEk6PcBt60A7Xqpe1E2cb7dpb0JSEShenuvc
J/95Iqy2z/xJmHj/xU9qmxSFMox8EvmGKtSYp3BBfglvmJa2AyHvlrLDFTcffPJ4
cIVgUNDfIHRgipaQlZfqty/NH1iwc2UPyg2jgl/pvyHELHonvpFN/yrgiVvEcUqq
6QESpKNq2+hBOLqZ2kBkPpW6oB07UdjEzeHrT7HcmxGWOb4n6CaQtX/0RIwTTUkl
wofcBLorXgZv8PYfnNFqwhnAnLdCxYNIceJwx5MUm1hGHVFrNQ9ph/9u4Tnpaw/1
iuJb/DzbfYkVCKVZqREH1PZ0gMLoFeBK6sk2Np6W3iF0hO0saaWU2ajjfy+TMw5Y
wIlm30kBr/ELcpzbdbsRTIRAaJFwnvAZ1PTJMC6BXPEuJvohkkBPtdBMBE2FqqEo
Mdnxsuyr1P2aqDpnbpA2uHrwcPtH7PgTBbqjpKhvViNMz7LCUKQlmzGk1FWb3SUp
p/yFhvutuoj62MOi58be46VESk6LqZSUTH6cIEWME44QSf0FpGyOG+tsAbWnr0Pc
nhkwpFmG+tzw2j7B3iZ/DT/66RihDbpcTrma3QECp9qwJ2Xjc8Z1tII7JgkqHIKb
iuwDK1QbtbeOvrgUBGV3uRHsCgXuZUoMkShMkAc9CiCP0mSquwmt/ke7GcdaFkqU
ReX3pSkkedY0FUm8Gq/PhGhWMdq0UqYMvNuCcNLAKQ1ncanIfD4UBGGttruignLm
uDgcngWL4Tp9CaT/LfbiLQG0YR3bUlqf0T9ImyhQc1qHblJY/ujtJTYqAvaAOXPr
IXTt5TqFUqSgwugRGZPNhcJs5QXwD/7HLU6ZlUIFRtfO46jKP+b2xF+RMn/0BiFQ
C4kaLi0Ie41bY4ycEaQiAgSjxO6ZV6y9GKJWt3wBpfQQEahtu7R4RzGYehIAwhwS
eiqs+Se1nOGqYLA6j9HGZGz+/nVXZS2i27shVYXtQJ8S8QP1vrp+dIaXSu6LZxeX
b+nxurB+WU5YXX6OJy/dHX7MpQy+l/nBHWXoyx0GRxEnVRPNumBK6yky4jtZk4OC
nJufnOPwCka7f3FebMY0wztJ1Qi5132nTFmphSd3SSku3O0yJyAeT0fPdRDl8rxD
Lo42Cqgab2QFbrdcSN7EiKzc2sgSNN5aTM7wRs0DKCv0TfteUtSMtgh8nPJ7c3/W
WGqNWSdz0+qdjH8j2O1G9Rlca9iBJ2UBzqp3sIfbdMyLOwJlFI1szWphUJn7LRAz
Z4da1nKxceCBmpTSUAxItNWQ6cQhxPiJ0mJMtjOXALEjg/6jYRsOuJH4/ucEGPsX
Y6dLHTURPehpi/lueVDu1dpcSJg2Ev+luE6TzAoUyPlOjTr/4wZczS3Ugg9SV0sM
sLgGr/w3TLJLpmzJ9G0eEtCrxqlznTqWEHt+4C8P83spCxgzdVqJcvBke6urORFI
uRFg/IWH4jQgaqIeMWylMMyST3kfm4mt/cUGEzF/Wx3Q4q3FEVTIz2GuwFIg+iik
+3wI5iAkSfXvXvdixXMJ2UJL/0PJ69swLFuZg7/5f1c2RwXINFVBFZi/TylaL7X7
7PVtnmhURYsWPXUmLdOY0SDnfGDmJeqKq5YxgJ2yGjQcssJCVfXiA+y2BjQITo8R
Ww0ShBLVxPd0CjzYBsLiwu80Mm//VBJERFkPtL2b47XaRUTDUuh/ol4uB2j5vhgc
rQ07bnvC/UvVER7t6b4pK5k/bTZJ3nS/DH66tkm6GDybFZ8BdDfvyV1JRT0kZx4h
b9PPnRZT2ySjNyTKNwixMy6z+Q6MPTXlXP7+4p82i3/879VQ1bmiZ6dH6Gj7GmdU
j0Q3+mLp+T+LQow6PhVBm2cN82F70rvieFi1SbJ4E7i1HDrKBPBIN4pJuAW+tCB5
AQeYr6j6DbXTdhA2eB3Wb9bmep9fNU+saqZJ6OlCAGB94b3Zv2V3lSSWHc4UijEp
SV1JP9iyb4ZOOZOSHOPBpEek4D6J1MkMWtgHDxiYyzOy30M4JMCZcfBJtePXvmhm
V5xzWYf+cclEO+SUktmi9rrtEu9mDZv2QMdNGD/eAeIMxbO52GhPuJYGYI2aPun+
GyephDUithtpMPo2Ct9cqmQM8Ly9FzUJ4qdGOAgt2FBlyc78blYFnI8jufV7kK7z
MLVt9LHN0SYj2OuXe5+D/1vZArjTN015NNpJbg+vXi07g7GS7i4g6AbpcDUoX5/u
C++SPwMM8KqKDSsIBeXmFP9FQsFZqpE//IcGeYNQYBZGEm5pLbTtpvkY0O9ZFpWa
+NCMF9lawMoL3VZjyVkUcY/NCy6KSi52dMr+zj907PyAdj2EibFMA2XKqyQRzu51
DB7AT9KFXowu/0ZYAovhTEwkoyfAMkJxJjHQuKAwF3oN9MzxjBcBIuEB/KXpt2Q7
dmVS2XPhApg2zAj7XU7nMa4gXTA3LDzuqbqrzRPUII3lQyQQ8ZMS+7rCNU8mo870
4WDCorrpXzMemsfpWvB1fSOnAh5942PVSRp4qM1DNF0td2LujcsRmrxwRndX1K+A
GkfFrjmzmoFYQIeifjTOdLDkMw+ikGCa+ZH8iGo6MtYHEbzo8t1obwaQI5rofjdw
wVZTeARLePiyV/TlzXAhNRQDdZDqVMYEoL5ti208e2C8myUDZ/o1pt+H69+6U+ZJ
vnRTjXf2PPq9aG8cyo8CfNlq0PHWb+n1tosdD8BHtNWU5Op0EYRlKNLDssgwLn3z
MflxgXZrJ/gd1HsBf4iulTa+o23sZg1khmWIFkAhd+H/argImwomOmpoNALGmox4
HPfEtzsgpt4tBFsmAJ9zrMVay2w127f4SMj0gDl7ZLJNVeoS7Ko5yKJUALLx3se7
3+Tlr7VXuzRTexAxMREFFeJdHJyEDFb8ASP0ZzynZ3XkzoSp43OFl9DGcgJ9bucf
OnGF5SzP7gMFEcisvB55Qdk+c4BsMtR7osaXefwxux8welpUWnpO+GNQn8SXqiI6
qT840FLo1rnvMIXCeq/BQcYq31klxUwmuAuGUx44uTTOurj9wBZl2IyI0TidkZ8S
3XbzK8GeT4/wR/l3Ww6SL8NJ51difdhrvRjBL7fnXb6v4/gJToVTOTt9iW+/NLL4
MSESwXUVtlFUV6wvojEdaypRMCIveIG3oIR0kAnohevKiaFdpKTYo3baFi1nz5O6
F3EKBY+zzkstNgAIq2DHS+gKgyFhMcMIhfybK4OFsNOAvs4o9OYeffd10hCyk6yq
15IXhjNfCTCEqByYNu6fMVJW0S4orF2p8rFy6OA88zIHfR6YtVnQgt/r9uL8whNL
SSTlcgT8S9CwVK0bfRN3OrW377m6n2uHDZQwFWTCOi44U1MwIswEUiUZwD0ALK/7
2sGUkwO45nYafaaxXTu00n6vN1pd89y40lCarGT6mr7N90sPQJ/3ASqJ6hRGd25z
Fp3KLF1bSYb+VQub4dCcNpmWAkVgjcNRV2nmuhjCMOIKbRYE0L279Bm939d8hfjh
rbRgjBrYvWwGCx1vainRtdU2PH40Nvq1TIL8u0i6hsNlskn/TVG3MSG+xde3a1GY
NadozFT48JUnZEj8UfegHCDU7QUn4ma10w9ndJvYUC1SHkI0TV/t5UMAIJg4Cooc
oXzDVythy7i9ptK03iKtPZ1AV8OIRKNXHf9ZrVVGhrYiJuwdpUTsR4XJgv1CQURA
x8OChdPlw8vikhK8n9IQGs0EI5aH/jXLBS6D7+9VxexoAvx+ZsFP7v42YU+JGAl6
9eBsZkY9RS6JEHUwQs2B1JC6087VCkfNtooSHJkyKwxj7PGc+V/HHmRaIWjDARzI
anEcJ2JV0BkZfJcMsB/1bZRC43BJx2aC2KqDT3l0ATprPnzZfTH4gO/ah5ZzYj+n
8Q/DZrAdKPtH/xFDQd2vl68DicreCq9WgvZX8ARkxUdZ0AAjb/jzYtz/7bNkUktj
mCI4u3KcPPOylx4+jzVWs6Q+d1l85eKR4dSQYVJlX31gO/3t7FPHs/eFLeYnfZSR
PMXdN6iTnCaV9Pe5mvxkp2b6wv33g8GrGo65L3gXNTWnbK/YgNEWaN1aDiYrAgwp
P0+zBHd1jh3QfHU8GoDPkB9Ez31ip5pALRYxIXYAvmJNGpkArEfxhpRjv12pH+vD
wI6OxmVPmi4MoXluflr4KS4l3jG1K3lm7XMthjRWCp8Lkw0Bm5GsrmW8BTYdaU4s
uPUFKgg+nJofmBCCeguK1aDz8wSonrTox98ArsE5szA14xSLD6svqGj3kgbKmOYf
eQsqsoDET2dl5RCkeEKxoiHewxmavh0ow1moOJQqFYe/HCP16+Hvb8RsICduzc/j
YSvMa8jl5U3mhdtt0TABpLytTiBesazYOx3l44LjVo1JLtj0eq/7J4LNVEDxmtHw
/O8rKaP3aXwJOJIDOUC9YB/TbomSdpBZZNtvccgXNwhvkiBQGCKegSW7DKuXk1Kj
Uc2ANTLhsg233+zvDzexnfrJe8qftIqXvFuFhA4gbr0AZv+/ifZwpZ6PO5+TYhA/
JdEXmxSmuO1GW+udOiTa7cQed+xfGFT7azRt6GFduXS444N1x9eOS0N0z8LYE4xv
xdY82inn7ij9stK8/eQe6nr26KaVLgmoZl25k/w9NfXDJHwoJoQhqslBACMRxhFU
Anq1pbKgrC1tDTg6jGPbCmXJeGzn0N13c6MUkkzzX26o8Hrf4NrcAAmWn4ghp0cU
fuw9KGL6jMR8xbVeuugUNzxuM6dKQ33PvWrxeYBeD9t9P4+Po4q1all2Jrq5YaXX
muf7J84v/EDsV2lmdo66rbv6y4QouPDyxUBLfnLmMW8YMqyxCKSdcuVQFkJH9zN9
vryTsfFtOIA6tkcn1pRTcTp+rBUzf8I9IO9s7Q8vOoxkZLS0JPmhXQNQF01zJ2zT
4b4glgbJBdjrPhMYyW80QKiDbfbNAwRH00mlFnXFR8vc0R69tqXInehhwjsFCMgY
jWuctpN8AipWotW6Oys6aQZ2+fz1XhZswXAIqltoi3ozonpzvnMs0pyfmvZlg72W
0NhM5+pYT3r9v+UdSSUs55bckyOqCzqCXFUHAajlJim+mvBrEZQNGeADIrdirM1n
YGOdbjTpFqK4dr8Mrmnwye1Jt1BJwYOTW+L9BRKNNPrq2XzMHKCVEik8x+QgkrIE
6+iQkLIUcti+R08Ir8br4nyJ+tPzUAnuU9UTXMC66uUXiMExRAQmFPsp4O/9u5xt
detjGw7XQmtWq8Oeq3EKejLKY+xzE/WhZ2K5zxwweMyx2DIXYoZRQFVRjJblhCSY
/ofWGb9d0sCOxLawTFqNljHzyBVE8ZImic12coMmlnrTfGcd2AmW4V727uVVdh/y
JBjjeta7A0bG/d+0/srd5D4+jRf9wwNpCq6WxGVYRLG5lAE6jAQLHniHaHTmMY/C
wc7vakrwEImpfLM9jeZMuhzAaKRK+caSNS0J+MFnp+jM6UIX1J9taWOxffrPHvrk
FtjLc1A7k1AuX8mMg/6FgPrAZd2knNTXZKVggH5FV1uXSvQD3mainBfGh0NF8Hy7
rH4sXxAsMpHNkDL53EbJciaDQCKu9a44beM4+uVoQVcMXVm5LyPAVnnN4qgApGhM
ystz7LyaTURmm3IQ7Dbg+i6uYoARIR8U8fKAo4/DuTn0IaghW9x4VU4dqORlp80q
mKfajHgUuCWQcKFSl5LBXGftMPRom7XFayNGO9W7j58Tdi4RxFyi++eOQTwRiF0r
X3fG2aHbJ02JFtDULFlxfE+goIyPcrugi52ClURJRCeGpx6s5Sat6pE5tvII/Jc5
t2yEbK9XYCij3Z6/MAFUDAr+aDduD62PV+HqqBH2BqRpY+1NyPAku1RD0J1kiNTo
gU6G7cYlZ3IjOGpb+JCbh1aUec+q27tvTfcXtH2960Q3gxp1CNFmnIS698y3zahL
EQfWqYyoqUsIFwGTKUpIjeTMujKT1hfYvb0lUmF17s0kqHnDZX1MXXmIzuWkreYK
oRad4rSzRIiriEz/6DMCDXXQ+0UfsBhqlvoLOdXzw/hgdD6S3/Yso4ekkj2qpP7W
EndQRWuFvCLfhz37FsRYrOQQFzdY6e1fCB5KxB4BqQOJLMQ3eETTzIvlStSw/FUD
Echu4MQ7Hj1yHm9QILWLD2GAHQMKlSH0KkqM7XGB2bd5RreqfDeQKRydTzb398VG
+suU9NM3xGttQymImJF7WvC68F4v7+oCm/J8JFeIl4oRlPfcl4EqyYpdZdwBMM9s
dO+ol0w50I+2/x+fNW5dt1ZiGT6Ssjs1GS2DpoZZV0XTVz6tckscnn3eQiLrWI2K
IGI5JGE+UBxzQr8w9A4ogLNb+Hf1v289Xl2Y8S+a5bPqQsVxtTOfHcSkOS8zZ3ux
xclrXz/Vhokr/T5GWyEq0ZQYSTwl8ruvMsELUYqjsvEH7ACw5ycKUmLJiOiABerP
M20CpGtAOZFUP84gU2wqxejTu+M1HaPLwW6TPYvkZlmOMRno8f12Z+ijWoqATOK+
2063qPmeNEqgzsQK+Qp+oJU84dEff5cU6hXLfz91qaojp8D1wzby0dYOJATXwziL
ZE/ijGKkwbutcWnbDAZkL8SXd1LxweRuU2Ngnx8sKIkdFeBw9HT4gqrIPiqqgj9L
CNceaWXNM+yaPebqzfWrEOUBAAKy38835RX0sHQejiqOOgI8xkW8rYHIPR9UXLbM
MrBOeGdeYSK6p5RP7cPF3kMNq7Z3fPqoXilvAwoOrnJdxag/Ro83C8OJYh7rpObu
Y6Gq66mNDWUnyfVXZxWUWIfzkFBF/jdhciUpHljloq7zuyg0WheOWoqUgTEI6hmy
iwd2tn8aV/ssY322sOJIIuN1QaRKhQXq6CEG5PAu9KYUUsFOW0WvTwWaqWnqKu0q
8JsZtksIjz4tChiaPo61PR/f+RHI8tLN+1wYHiiWRJv27wWO60oOILiS0lE1yIKM
a5LcBE3ECKG0bzB5DDPTGO0XO/SfpgSFcV4jLB5QEGdJ1Ic45dQK4kWVymqLmSmD
TLjZXXE05ofyeOI0JIhwFelpXHznFYDQOI/6TSSLvtq/pQ9JoR5WFOSX6WdnwzsK
sMhFVQTXIhLt5ylaeL//ecdOAOEse5BjyTgeHU5RVQUPWqyCze8sqHnb6jrSl5m3
yXSAWs/JB+RYkoYcEF4tTN6IOIvgiLkHI4uix7eJN0ztjCBBj3N9uBpo47DdGENJ
wUWoQRfVx3NqeFN9WF+a4PcwMuzVx7r6HGbWo71gA8gqj9ZrHZWaDE+OpmPeW7Eo
ShUDL/peMiD3pbmjsxZ5mnqqvtIvzgTtKatv0Asu2hHnKNtOObhHw/h64UC62Z7S
3+x1mXjO3mCA2zcph+lw1b+RSp1h4ef7qkPoF5AKyjunrwEPtOTkEnweetWsQ2Hy
SOrBMLiGaEenCJDOV9VWx2gfNZqttCJe8OStG8MAtPJ961uUImX7mr7F0tb2T3Jx
ODyb+dMLUYlVS3qKCmZQ6WJ9pN9cXVXWEmLWYkZH7eUqYlX5Hacvv/nfw/hSsmu2
IFre8AdKCSv6pR+qvjDqPCQTMzoHI1379oRlZ2816Dx0LMvdLcSH4QrmuTDLqLSA
6ehi4VyFrV2VOJuDERCOKljE7x7KCpyHY6CDFNGkOkiUBNMHlcPGWDBkXp4+b8MO
JfN9j1lGe0P2aUVoNQFnfSCD7OLpCVdNUEQ736iJqzpQ3zU9zk2jEyOO6goEoQxq
L867YJT+lS2SlqH8ANSqG0j5kxlDliulK40vtesx/kXkBkc75qXG7FdzBly4GK5o
PQXuG2n3liT3CPH3oX2kt/Z4fc96Esby45SyoynFoZ2UB56gosJfTN8ciTDJcmtd
GBTBOk7R6h7rldjc+XIV8SeFNpceDKzvhntpR+bA4d2G/494f6tEPTwFx3KjD+Qq
9Oo7oUsHZclBQgSOk7dpYyiJtvEdMcbkpp6kDx7yfCHP/Zy2V320OQ7fB8RJO2jQ
yVZGrImLvPH3p4seELdFoaO3vwPz0Qm3CelfW/T3ZWYQh0bjtg2G1Y4e4rSR08xx
nHQHnhNDp+eRcLc5JjjaixNgDbpp+JvqmPH9fpTqa9vB6Nu34cJ5qTUo/PkkAqki
X48R9oVfKm6Uc0Nxcb5Btq2t9qqPGaJ2kZL4Y1OV2yoSzPa4aGHt+zIVfffgku2r
x4SHMrdC8ocSbiZOMq4yqgHHuAvGCOf8h2RmuMbtNMiyF4Yb2nrtI1Ll/StmpyoJ
by2TeFT8vcj6cC5Ts6sY8oF/P3XIGhjy3EXGrvCiTHXfWbzodaG9/gMZrFC+jztx
qLSEhSMb9Sia8uTVFYe19uOyz1e6fDzH2xcdBc4Zzfs7fsfrgZlD3CC1hGYD84ET
ma+Frr/GLknBJuk3+1sHukGBUJuUCM3bFKDATF6pUNRgoIjDpue+Ms67KkBhiF5O
kYROcrmnIHNQ2RGn0LxpVoC4/tZ82tgBSY3Ne7yFO9vopSNpFbn7+N7TEIAfFRy0
S8MeDDRyaDgl4gq+ONIGR6r6AIpd/119tf9UTHnLvA48CuJZwE+aGbqGWvnJSpR5
RIDnFKTbmEHJG99vCHSIr3fjjqKvBjIRauxwWRtN7DuM6yxHD7wDDF8t37cJOHbk
HxvGaoU0h+cVqUuUjnEAc97ufIMlcV5QpKGMAylz9paIwb9nS3ZNlNXfIX17pBQa
22sFGXPUsJvzzypmbxtEREgOPeoz7X5ZDV+DS9xSJFRhZbeRMoJIr5/XXb7a9jpL
QPe/7+/UCRxpxG6FMOMQn62w3FpNjq7rGCOEzkhwSlfp3McsATfgcxFPH/Y0TOWA
Q4gpiV0b7EG5yjuewiA4WpYKjj+Kdm/wK0KpVAXXAyQlbJE0R7+5LuWQ8wFKF+08
NaQXqVZA7WL3IQoceSCav3gxv0etyRSL+165Ig8kmrpvp9Wz70e9z3Ov8Q2DZ968
FXEizzPxAzdGIR9EmFTGRp5hceXpC1rLJVvmsDosp2++a+hkR1dUQJgYw0alrNRU
2HQoisHp2gdAE2hwD+b5M/2y3f9ltkxT5B+W9xPxPjM4Q6jLNDlCASJ66xLMZXSE
ofcoHh7bxRHbDDNiis6i0VwiT17+2RhtuhsJHZze8ClJlFgVabaJHiowbagtW+NW
WpqoFyMqWT6kCfJO8Mw9Zj6SAHqo3LiLmVqOa3M3R+MuvpGxLLXsgY+uuHwhJPxy
8qRbGaGTBdVon4Pn7H1+awHYy47PcsAfVkV/XoisBFF+taKGSiS9HKTkA90EUCqX
5INgpiAOj128V+Ui6X8hTJhyiAQRJzea2qXNKeBN38T/6HyXOlf+K1cCtPtFO/bG
gU0Fk26/rJrrMG6FoHGoethT+Pucu274QklbURYxRsUCOitXpFJ+NT8cWh0UVrg/
THnZ7RGSReqNITOxmYSnW+34an8OKR03qAlUz5ND6Q7gAp21zGwKMeRXtOpgWU40
2uVPBzYmsovousNm7tshE55oH2emc+Y8rQqnFdq9pYDCbFJ/s88/IrUEPiPhVCW9
OwxfFv5bGh6WT4dzmLaWo8ajn9wcQBL8gAuHpXj96HGP09dVlVt4fq7UHrFgQDxw
oCAHb1ZyFWvoxrquPOeZgSWL4Qs7QDjywsbc/I8aFhYuQRDlkpDm9HEOTsv/kQFu
ygmDkjZE8FuC6R7+c5LHRUAgAU5xaeRsHrMI40rmRttc1kv7tYBfL7N81Fg/QrWo
NGAJBJEjaTVcErpwB+KFdXv8attYVUmx6/USDmXv5FGR/nfuaWd4NqWsvw1qnIC/
ULAsNkg8mC14uhTlYOvAC9MVmF4ZHs7hA1jxMAFmhbCeWFe48d13LnvhjnwW9wO+
Czi2Arvc+tQsyXLMOgPkwagxOhaFuSR3hNoyHgE2uPlUYGERcVehO2tBp9hZ0fWo
nWUaf3P2/0FyV6QnmOMNkGHOtGoWHExD4Ub5HkrTKYxrp5+bSPO3Aj1W44t3WWJn
98EfKgFVre+5W6B96P+Qp1y7RShfWgrI9QO06PRA+d3nyC8G8W2f1hpfio8I77rv
LPU7KRGjR8E6ylIn0JasKjeN5R5Dys7EA4WmDm2vbTyT/UE81Z707uc8lKih56C7
r4Hp8wKmHv5rXgxrvHNsWR1Ijn/dHnXifq3Wvp68BbFNWhkFkmi+YCywe17Az7YA
jj26CskC8hEGOus7yJB6xk6gJOiJ0E3NW7UO0WpUDZXslGMkUBemVsIiAKGQz3Pw
A0NAp/W+Zeu2ROJ1y8Hsr2vsXtjKiFTh/o2OD0jj9bC8ycMQtxBJL4/blvJC5hXc
rYnMet4/Sryg7y5tGQbfXbr3oE2ZmXzcV5ZIpaRsUp0og6a8EOcqcZIzLMhwqKFq
MnwF/XIJAlkyJaXc6uegIa/AeWHohid2UJ0miNL2FoCbGM5iANN+g0fhEFeGbVnP
RiXu8EvAfb4Cef6Xkr9lCWMy1WRvmdZDbJ/0qytHT1eTJ3rt2WkCCND49dp4H5cW
YRv1DazGXVOGWD1CT8BQ+ys0ACv41s9a3UNJDpPdBeaLYnDdV8APoz47bWtmQrRT
ERu5NnipfrIlBoQaa8kWOKfeztxTdTT1bCTb3VNqgTSHuxSZH9ELWq+dcVUrr3l4
qFITbHmP7hFdRkT0RSgFbQlT09cRcHXy6RPz7hHJJzGZws29pBtmhpCBMkBwLv/o
oikFosx5KLpPsKb6EQLl+LNIHHQ9mW1JT+IWvStg8hqCWYqLzmLcSIkttaNPps7g
KmPoVJRe3En4ewRrHCAidBEPxRDdSlznaR+ZsIXIA7Oj47gmn36yNJwXQiNnMCdr
dM3hP/2SVbnBIeFBU9OZsukmE7XAXkApuYkCXi0sodrl2v1KZR7O1AYmuDfjP1wZ
uPWSD6/SG9NlsyNo04jX6yqA9NI9NH81jd0MtqG0CJfF6xOT5vS5AWfPgNFgrxmW
RMNqw9b5/y0X+vCgUr73KKAAdSbvsYi+rcHXEfLqopXL86YnuG7n3mXzAae3I2GW
4bbpGyZbuAoJlyaP+8VYXg8l/YKi8shBlIZOCiPBZEuXk26yTYJheI81QoGkodLt
jmyamBf1xOL1opTl2ul4qpt1Vs2IhPfc60K5dh1J6b8UJghS3ULp4uMcDyySH4EG
ICBO/asQR8Zn3rFjg3qZC2A6RxDjIjEzsEXRmIPs7BnujzeyJHPATiX28+87XJ9t
TiVwfD/nUUxGsoAfG5n4vY70ARrZskXvUPNnqGtgZ93hgEa74KUXeiGlhcOIdkzp
bggK4gzyFPeEvr0GiP8nqr+tWkARlnJw2PF67FL6JJ5fAEQQMpkrISWSLsxI5lgT
1usTm5LXnjfpS1hZiWM1GvmWFGwoZ0LnO/igs0OUSboYTMvf5lAO7myWOBdp+pDD
wsETOIuAa642sWQk8VXyj+zwvOR5iJx3nH9tqRqW0X1CSeBs+KOQfOZkEUg7aGzS
cVdlKFmRUIv0SCCE3J+/YVoNiGv3h91rQHWODQMupGoHk+p12UaZDqLMfHZ2bhaJ
4l1Z7jFznDTtE/fQPyPMjsOHwFM0W6xrGkfu66U7Oc7BOB8ZiuhY6u4uJVseggg7
YUgpakwz8ZUwgZPtjhP6Mj/DzsuyOo2T+0h/kjCYftETeGwcs/SwzvL8JUVER3pg
+gSW3Clg8OZJI3jrUjdFeqBh/gzVlkb1MR4IEB1ZbopOwcC4YQjZ+Y0IhOXyDKqF
b9OtJs6Lc5c73OLZsgdWULpE7OTb2tY0rOaMHWjvJ3dVT94vRS3FzDibdpkNwq2z
uns4nF4U+9KXslMTi0jlAX44APgLQx/gY27ru6nW18XJQjpCl6JesJiJL8PB0r67
BTL4LBBiLEKeplwWSqL3oVhx636RmNxiS6uEKIKnhWWpyIoKgHg22Y0V7VXIAcrL
0SjYrB1TtXBQc0pDFcHskIzE1wjmeS/V1E37Sq2q5a+tIIwNtZ00sEN+7/r2HomH
xcCnOe8WQdlEytD6VLPemdZZH/tMTJNM7QxYH/Do3x4ZF5BeLI81Qzaral8rsxvW
eGTU0PBOwrZ3GmjdvSh9bd6UWiQz3Lcv6dzCaiZI8EnobmdMYU/YcRHIV5+YTmey
V44osP0rGyXiIAbgy0a1Sd1Rss+tlbyzOXaVBJfXVa3hxwCN7/1jWtIU6ytl3EeC
y3h/FH6jmxvavaECDQfSYqMt/G3/t7OQBGgGXOSFpArA8nC3oFm3KoaXa2H39tV0
xsmBdcuGb4TUqR3njSs7cJLHyPwHoi6ltWyfzhtE0iDOg3yzGhscZ/0rmY/ViAm3
9twM94xNYRPQTsqEUYLxo6waml2BZd1pXikBOmWuiznv0YuJ+ySIWoi9c1ZgutY/
TYDTvNjHrKTmQsCRaG5QLkx+M/A3AD97UoWT8alKLx5hQ+2R9Zal2+5WZ+xRnK6k
2Lfg8o7662l2s0ProoBAoQeBEf8NVnJpNLRwyqFJxzUZVXY6sVaVYgvz0FaXNhWi
+vSndlB5XE07jR1AOoYsiZaG1MLVb4TjJp+btBClsy3YaLibSKzzOh1iHxIFwc48
YZAIAIyK6OIHP5uDY05Di/IrzI+EmKmLDSBzLndc52D0ob1Wc9ICg+NoZOMi/W0h
M3waJOgiIRy6sXk6MUx40iNhTrDj7hzqbB44qUGWMfXoIXkjXqLCpk9+s8x4O/tH
cmrc4ccK5pYo+2TmfQYboevGdsNWM8F1dc5snGPaGPqQkdoc78SHyAIwS+dEYfJA
0mo377upJs1rXGQg8tO/6JNzFoBK9JynQM+2RQirl3DXShlKtrdUFysZ5qBZZ6yZ
p9B3SWBE3O3TQMPnDDiw7g45p/P3NK3keWXK+1qcyRCAP2zMLZrbqJpga0uhVCuE
flyel1BfdLyTKzkonzE3zP10eO52QBagncWs2qwZtVmTU+/BEQcNwZ2EnYryzR40
HBq7hgLIKZmDhm3ajho28AIwpRo43GOCMkovQjr8cit/RtEIAgwMmG54IAOt5hkv
rNfb8O6FjLZ9B2PVbFQVi8VAQj+rJfHWvXBzQoscoatSFV2MNXwYB5Rg5K824bpL
amgIWaqnQOg1u/FnuklJmdgyvf7P1I/MB+b8ED83VH8Sm+3yXTQhkF4M+d7DnAOd
lLFmtrLMLkgLe9zd09yc32mSs7JsfqIX3sB/KR4AxcQxph9U5LDHUXbEToK0TJ1Y
iB8TMT1dAgNoPO++409SHQG9xJP48KJKw6ury5pin1NjwESJWRo9rdSFUpkmq8ef
fvL41xF+Sk4fFqkFcluoVwOCnbnSAA6zAgyoT/IGfpkoQp64Vw119wsU5C/B+jtO
6c4GKRPKrhqg1GNiPwhqsWbu3Kq8tDaXvQ0AXWKMhG5Tzryn7J1kQ3DPJ5upJW1v
TZ1s0meMQJ/DpucYFZ61RW/MQ/zhH2PczP0ZOyxH9xRyhwVDZf4knLlvCDlL2ZOp
STeIA6O991FhX0h0FzGR/xqKTZ3Qq3XkHSo9Y/stxawTn0+rhMv/b2pBvfcd1ySJ
GHWGyOI5TloXUaUz6+pvBE+5d+ByCTQsd8ApMe0U8LTnWt65sDsjtR2id88ivDeD
RjB9c3hCiNFiynuojD6ySlMncVADLDzPTkO87L5Grpxr7v8KjnsOL/kJyaMuR8bf
cEi8NPpU6gM8DvsEGCTGgEp4dfKm9G2Rj2svtv1wlrmj5UyNtrquLZH/F/dsxtWi
CcpmP9QMZ7lPAdCESQC9fMX1yD+/cX4kjOHrXx8SdtRcfkguFtO27a5cimSkwp38
rY98Ws52jYIBTlHKfKxQp2V2GqohzU+gC2FYEEXKXWSBFsO/cvTR7puAzlztfbVI
cZ+ECtHDl/lVBN90C2UESZ9e6/1Bv3X+fyUP8JvVJv/5Wi1S/EYOfRWpI2uL4Aga
87TckiCK2TgtknDJTIEMBjBAgHbT4OjcTYkwZavlx428pf6oA4dx/3P71tkmXMH8
pL0N6ZuO3XHKMf6gED7BmC2Vle5P7cKRzuICs2OkS2UIuUK7BHOaqzTYnfrKEpQZ
ubhiNw+CFvrSLSxZKEJMvGEAqcNnCDrWRvXEeY6cjYNBcz+RqEMECUcxqahMFVqQ
S8KZH0xbxlLBWphdVBZdngciOdroq3GUH/sqq90VgEzeCYTF2dcaRt32o/4uqU2q
U/0Igw8VuvLRh65M2/EYNXM6dZS7P67Bw1lTGlOFoawPa2MwW/R1AFn83khemneM
1XR7I/564uFvKBC3XmJTtCBTQdgboSvoP87a8p3BiYW8THiZ0A0HmNMaz7LrN7hP
aasMzdhb7MHIJmGkuH2w3Ej/u9ruXKVJp1DMFlE3Ic+2uurEKjBqISLcqoGNEVG4
hDWzlWVH4fBRIhI8WW9udmJgxM1f+YXF50KvwPYBu7m3cyM+r2F5mINKDjA01E9a
Eq81wGf2yp3pFrGOJySi8MD2vJIRbnmEkkuzasCgcWm74Ma/SJRkjohwEU1iAZ8J
I+2uCV6ew2TLOdxHY0wXzF7WOZ/MRWEVBCklBztZQRVdZgw4XDRNPa7iA7cwFzG1
LvmZHNs0O6rCPUGuqyjXBId3K2c3xK7c+11pd6BBP5JxubmppalaokwBIcdU4Igw
0tplY1JhA2YplEhCVRiynF7vxYLuf4YwxnCBG69dVwi82RSChXP8yt2zQCilmH6c
qW4to0964wrrnNOLpZEMU2jMJZcxUgpr1XoLWboLkS1em2Dhn5Xzfw2/nodIdHbr
C4LjSS5ryVYtXSk9l+drthtRgmDoazLxM77z9T0hbDsVnYhsfSIVSaFvKTZp4lAU
03dhPcxnobJ5pp2PjuBPLHp65q7dydFeLwkEw4uuAWPJeNRLWJEBdODumHr7Vj8N
xgxOo+oN27mZ62vSbfxdZVytOIjTUa3yWODzJQq3BJQgeHsh7K8/bIcuUbFqjeOx
+UkpvuqtxzDuZRHa3sgynjsai3cwq0lwI2tcTF+yQgt0RcNiBvNLNWr9mN+ZnmqP
62jgpxhRhWMTa33qlRF2DWHuTaMUFcBE1hxd8J6sj6kK/SOrCiRmUN9nHIB1EXuf
8r5Jh4kR/CUIBdc9/EeAoz8YDJqGUIimhwIm9j0CLD+hwCeTeZW65XxrkwdrnOfY
vSk2Uul1FfS/djElpC+NaITiKegDxzOE9jzEM0yw/TtUdwfIt7VgpNbRMkqCQC1N
jMjtw4BJd8jiZKy2FueBwkLiy5Cu7yzl/faEh7KUxH55CMr4Dlmqf4WNX4LqsBHy
nNeYfk/qOopSTkv3hB4h3eClTQ5MlfVj7uhIgLFrx+eDpc2QCJM0sZ/chAgWQ+Gt
C2GDYTiangYalYmS9VSKWgjrOFDRSpFBxdw0nFDH2cgM0cauQT/AEqLPAq2b8Ujm
MoMYusJMiewSTOsnHfdz5S/9eomZTJ3EkARJWqyjyUDhc36KxsAESlqvAxGy83Ta
fq9qPNZx/DAK99Xl5ntqE8CQ3DeREU489Vfu0Xe8Y2f7JXNS6ExSMJUA+HM1nwk0
57Sd4RfxnYgkPHsCVHSYb8ffzfWkj/uug9t3kLN140lklMUSB3SsQSOdP/tZ1m9B
jIj4EjL4IMhqymoQNwEhs4+vDbmQ2FyePNcxXjWM03GrFCAz+u3uGTc7aQhfvAlh
D40i26BW8iX/nl2v79AIkQ6VNNTzLsbmvPHXAAYF5jka5ikia5t0hVYeK/gvl5sD
croUG23aZBxIg+Jkd9gd8wvNjs62CuQLmtrnzv4NP8HV5/zAlMX8RtmzrGVTcgvO
hkMJl1pMjNtIbJ8UumbJTjRnccYmNnf68R7qddxgY7IFVWaJYNf0h5Ukn7ujhXI0
Mt97iuFj9xmOJp2PerQTpoq2U7YwJJ9hGOtNdgNGQfopfrZcSzvC5GF0HVC20Fsb
nzGjMid41EuveGJlVdJhh0jc/NxH/uVQQ/EIwNM/4BmFl5rASZIyIHbzWKDPKV8Y
GSAds6XjsWtwugbqFrSiNxr8mwYf1AkBfm7p/NoDcSWzgoB32//Ezbq6426+f9JR
lHPU9o1ACgWx9Z33eYHDGLzzpKXz3njjHNyU3nNYmKnLNr6W88BxqgVaKhMZi3z9
JCscKC4AWD/MhXfBQpPHcKzNyth7LsGGnRjlMdF9yyXOjiyOYpOSGloyf+Ex1w7i
HOW2l0IA3QJz90DabWol68t3gOPKJFSD3ZYj8Hq0iB81MIiKCfciiAZ699uP3S8/
obFo8nkuupx1rVUoukNzBLfIM/q4a6y+XDtrWe0IUxMMERwzw5AVv9LkIYPHTlhN
kAJ8OEmyDhxbBASqLV1oy8bQW7AMIM/3xqqcSUyYJqSLFM1QdZv81jqgXHq4KHXm
jUou+l0xMC3a1kjrFY8Kl/IixMuhFvfbH4+aFp6VHRyFLo55V6jXOBckeyv0x3DP
S03pFc6HPZ7Q6YV40j5CFXL1yw7H/q0xcOOeszhkJGtr1pbefxsrsarWg/Ds2mL6
yd9rVpuNawqFmzL0VE2oxRldt8aB8KT/HSaEdEfix+Cm4fYQOgrLYEx5OVJUdCRL
tvIl1NW6iz9XI89J9krqwS/lqhXIt1sXuhALUeZMQsd7bvxgXvLR0VTYlZbBDRmV
LyLg7KDO6/Kni7pngXsGrwRevlMwasaGxXgqrmgNm2IFtgoWK6FO5MlGn8Xd3b1u
8lxntL5dIivp/gdF1zeRvjYr5Arm1p4mM5vwKQQkxfkUPEsyIQWjetxw9DEULNyv
Sw4rL9nW+lxsj4vUI7lHcooXquaTY/u/JFqRMUMbYP5v8d7xU2q3Z6qgsi/KE48I
aqe32XgRjciNKy8x5fDTKv4nbBI/502SfmFj8IYOBm8jVMYlyELGX/vZYNJcF0v7
ilIRptScSqK5IVWZgmW7s/OeiqwyafokoW+nnJ1uQa+RqdWT1oqzukp4QFeDtGbb
lXTs+doGl2FV1CgjLslHR85uHVuy+zM9ZmwLfbh6MHMzG7xxLmU2iwp+i7Ry86Ru
IMWjCqbEAFq+CRdu9CMIp/h5m4DRPy71ncDVEIafAlf1H4xhWcjYWFdqc4QhrroT
d2YJimL1Yx/0yOR5RziX5Dqxenp17rLx8NexInm3NVIlKANEibWhtZMUrQR0GLPx
GGmJara8mVBabdI/1XvatnuRHcJUZHA+437BTeR4cxDbCWLi5+hHQ82hchjGxBeL
nWUTHwlEapA0I/0PEx4BVtsoebFSOO3kMQFFXwLmurtbuOJx3iFpdJ87kltzJnBk
D98wBqSYRXeYrc71aXoLzoqs2z7fxAU/k27Wk6vLUALxdx3h1Zq7i1tW3qzNqLCD
lIepKnbPXnnbqn83nBmIB/Qo/Cs+FFFu889+IQmuBGi+TJvtSzWehlcjA346g/0k
gXYRVMuhFKhoBgcHpUt+CXEWcNEiHQrrO8lK7hLZQkj/pAx6YpInEIhAYOohI2AT
kpI7DlCWLOrr9RGKOEypYT3gJyoc989STNdB8XXgd4lJVmly7/DNJVEMDkVeXHG7
z5W5sT0F4I4M0D+9v3TK/2GU/RNjyVVtqxw778OUFo7IYSiQ3WeQTVxWcmrddosC
eKHQ+z8/SXjHMcZM8B3X8Fr5qB2K3PHIb9WEEF5IYsNmVfUUieh3d9pZxtu6ay7o
S7S+Oin7f1+CdML5an3U0OkLAVHJdVfg5UXP2/WwSWL8LEYTQb8Dd8i2Ld6bmq7c
znILrTb9JB33kGucxs3nTfbu3a36vVHC5yJDOck2GRVJkeqL4xks45TemBrwjgeN
FFFs/+s1W2N1j3c9770pQBtZxVCmOLyqRN6qGQ45OG30V83guiv+Z3S+zzNP98OV
EL8GL/Ri12qKpw2NSwjcNHkBofW0yd6j0uDLNDF5B/127uECiTp+5lI618dPFbb9
dKDSwwqlhju8zaUms0chh+uWA5mkSqXu5pABds0/5zPEnAQVbBc5nZOVmiwTK/v0
VKdvMziHm5jXFB0YsggAl/XGwdMbrCdSLeNAIElULxaaOqBL7KaCMxTi/AJb9Qfj
MIqpilRd7y6PJCshhyDHLWMCb0CXOkvMyDKE1yFjjbOeboQAhOub+2mS2jfGNZ/L
gsYys1JFzOhEYeigqQUute0KmOeBuXE1jPtvVl3ThyQG/C1K5EqDhK4lsMqL62yF
LdSolyyM9WQsIibCKRgK9NnoGpaqe6+T3XZf34z273dDocDEysoNGYe//nKcXnOW
/61UhttBZlCIsu6pzgDIVoc123zauf8piFclILV1/HX22G0aDHEi/XUjNOKa7YCK
rVphYsS4t/PPB8HBodS6y54ulU/qLZ39OOuZlqZZD5iqBwxSYg6TaUEaYVyMrSgf
duI7SRwbH02RiE9uCHg9QIFSqqV/JBsfb9m9vbda13Nz9l1gaAKz3OOuNNU6BnM+
q5O4tyWZOonVpRd/gLH3kEZXkGrF2nKmzbzjIS+eyrjwUwQlKmfot+PBh7AgqHOB
24cqybuTEn7yDguxqucRN0EHRtz/CyjY8jjK2tSksa/TooBJ/C4+zVWiK0fc0LxW
aeyxAxKSaFPhrZ8ADXrsrN3fhOiyf4OsCta72HG0YhEJVNh4xgk0TVFHT43/n1rg
q+i2zFVNLPOThD2Tf7uHbnADa6gl/95GKKkvSOdG28v1heO7skXK2G0PxZ2jsNQP
ThwHqPTCuFGRRF6T4wrGON12fg/W3l7m5pLg+8AK2gxumqU9yneS1f8MTh8Vk3AZ
J2gUHxc09RZhRMmmvT9S4clOg97PwDY57C1eNQzLBdCbfW2BTvdGERJH963TulNp
k+BwxGZchjVWtZCMtMa3j5iaZmBKAlwMwS2RzeSe1PiySXYcwAAYyYxqkGBX4jJP
HWXPBIT9cXH5ddtd8oFSNPYKim/2YNDb260RSkMZP17R2633rxNB1z2Z9W+iBXJC
V22yw5/MX3YbT33Z5t/gCQ8NunRCx75MSjuuMoVCx2/yFmB1we5Ii4Q0Xg1cXLxU
MG21ItTkpValQb06LHEvnsvMyr4mvR6YpDz/FEvMon0wonW1lMzrJe9aX1qxp/uR
UyGVPgIl/1HH9Z5LMLjJrL3AsNmGmebynXu7qwvJWAKayxCtVkfUiWoyx/T5lIAk
bZmxGh48eLcqzUSYOvYDh3cugpqOkH3+OGLXPX0Jo8OiMlhp8lM3yqs6C2/m5XMU
x20as5H3uDT9kRtLelFq6s3Vc1vpg3ih16+gIXmaz88DcRHNKZRX2vMxsC48dN6U
2rmMQvGxlsr/hqcR/uJmf7IvUy0Y9N0yV+WjKcW/00GEoAP0JdqCTcAmqTAcrXOd
jvAonSk3aQFhSB5iYTjaG+bwcG8qPJKHohwoyO+d3mjdcurj1lFlCdVQ+sAVIjMb
4t+AGfidSawVAY+Ancp0VY11V07wO9fiU6MgoABdbxUcrTPvY1fFwQvV5RZj/wfQ
2g6JG5yW1VVYxoHJiJpUmgHNvaaWhWPlyRfeo7X+QapGLNSV3cMVAMScO7M74Ke8
HfuIXtYXBNhJGTVBlq5LRYRmYdyKoRhE1zPhlQ69b7Fo5dPh9QjrdHZ0zH1nRDAZ
IZYgcFj8kW0bnfO+8SKWm2jYSdAQrd2UHdhIYdQ9B8H9rIbl3GHJIj+W6yrDXlo0
8MMGppxleKemluvewqAB0XKEWmapJD3BoKVqcG2oIeylOiOjZeHbsnUDGXYch2g8
ZI/z6UMsxkhpVy31ZjeJunmxU60KGn7pc+biK3GK+PW3lX2pIcpzBhjH5ODkkXUU
nxEmIamLmVGkmLbwfj9wxYnwGIbGqLnTrMQz7jgZGI7LV1uVccEoEReok0GHZSQg
WfyZd7Pme+MobIE2VF/GslS/laqj1ePFAsDgt6skyVSosrEKtoeSG0u2krGOantH
5yNio8hX3cmPs4UxPb+1zFRQDrkRctvVUu8Oc3/Wh8HhD72kWgwLcrIyAURJS9uH
VvRsHpV8oBt7BIciPgpOexUwy+ifrKMyI8cIDrEkAm/BgKBlA700MDaBY3n8A3PH
ITQiK1tJtVWiqrApqwKnRzt6htcOzIOpvyDAhD2JULgjmn4eWPZx3XJ4F8oay0YK
FxHJGECuIxT5lgn/6X2Ceb3x+xC1KqnL6vZ70OWg0H99yw+LEzgZR06x5JVNLMuP
CE2XtKjrfRudzxcvneFyQ4qH5DWhkT7xCGI3L/34qWyLofUW0Qdw+HvBqAYON/ul
2Hpe67DQlxia8hKSceADrNL37bXAsuqUq2GVlCdpDefAgmFpSGiRBWqNVrpNMBdM
EDTGZtHves69VXmSp/dgVlvozstJ5LNRvApfr+xG+ULksRoLTaleOJ5BTnoVXP3P
j+sGF05EU3XL9dwW/PBsK4LkDrM+BAl6PoHGI3800Lk/RTDqATmIC+2wU75jc3rO
GX6ntpAx6EkngD7rJdtygjvlSyKItExw5fDBWDqDjNrQ3xyWBjcxYOZ2uT3FlzfC
13Ax52QQSoIsDhYt8yEFw8N4ZQkwFZ37FpQPgeSRRhyuJZi+vy0vNSIvK2c3Idr2
yBAxfz2eYTCcyP9v4DDZUvOmZ6MD/01L0L4kwHLJlmxVTx1TQhxZZ4p4+X1C+7cv
yF8Ehi7ul6dEJsJFPRpyh3bUmeUIVmLXuUsj47qzwJCtKo84F4s6OJpgzDGn8VTu
h0b1vAw5lJqphiFrq0ORrtaMCmzsiHYuJ0yUb6Z72K83CBJ0tdjX51IO5WbFblpa
34nbom0pCR/V2Fk9238Ch6f3QRP95eE2bki/Sh9CZUUqAuuu0YNG5veD/poRwF5E
u7ca7wcUmfuPvHKWcTcvwoFmt0ELbzC2W0od5yoaAHSiKWuJ8sWJtLCIiOma8wxZ
uv/wvYK8SvTok3pOZyLt1EDjWEUfI4ZEZgMW/VchtaZT752x1wmYhYgYbAyhG1kT
1ywhU/ZJCc0Ej4VitCkgSFBzCl5q8z2m3i5aMsKZXs2sVf9Co9NxU9tvNizxeaYS
AyiDAmEVNI9AoLtrGCyuWzjHxE4UEsiYEyUzHhvcBwq6Ybrf4Z85i5pMyNMGuHBG
Ygve8bNDZ+slnxKCVptuJKFUBlEq0AT83IUm+sGmG6SoBZ3kBIXnPRduu9URYNd4
EUC+rL4n5ejFgkUx1F0KVpZMgVDZ/mZwVxAD9zEfTq+8CWMcKX8T8EBEJYBp7btv
SyjIOzTDUhN6humtDW72DDTH2vEfFfSm9TE1i6GvfddbGqqEDgpiGnGFpaGJPzu7
DNy6WK3w7yJmRXtjg6cpDo+Ox4n0IP5dQzbsQkp7J1pgTZRSFRGJVWs7hC4RcnOA
UwKXQZ09saj+S4NN8TofT9ef11X/2bDx9L1rFXmlShjkLY2J2vslgOtA0nRgTk3A
Q9EmRL8h8ijcIBM/krbwk3oAUKIewcM6R6BcqSohUrpJMQGjSXFyBRRr5Dp/i1Aq
AxEdsM/pXjL0f0a9LAH2ui1lpZhmuFmRbJp/zWUMeqBuw14IlwAH2djpLF4/mHSA
uUpg42Xb5irU7ou0wuauulE5gz0zj0Vhvc2rfY5pb5ku6MJ09sNe2gxYYafc9jWG
qBuocbj1M54syfszazrpG6t/q+YHJ2YuvuKsi3mqg6G9DCvwreel2JtJ+6b/+0fE
4Q6g73U7YDWpXRVgDSLqD5tsbQxLlYRYFxBTOrmOkjN8vzXwtui5DV4iK0huPXb9
RbeAinbgqzje3o3Rq5CpASKvxarue3EeEwi27FkFMOAUTmOgtpsrv9kl0dw2ueik
U63uRrNeCXeg9lCcxcRCCKjfK0SdGyT/3GzwVRNUmne4YY3MfzzmV7vGVJnzpHdb
k4f3dh0YW/yM1CVNQWVFYyMahQ4TW7ACtK4i5Tx9GPfBdqDSiWa6mv6IH9MkACVZ
BxFoGEAVwQsN1PuAblIYmOXPKYIwZ4cUEmynyyKW4Jm5bay+gY6UO5Fxf8xI4pCP
EC47sOUi4sXSXFjxobTe+rowv6h8BZkmXDli2rQXBauZL97ti7wKYhBL3PpXVrzJ
Zcj8DQ8mYd/k19TgLK98c2ihMCE6Jhs9EWXjGsJNalIi+B505wiMsmdRZ+bvpLwr
t4Segh8BkaSym6gUuX1lGwXX001YJCSruZCUeK+e7lTKP+K8yU0rvAjHbpzfYSgM
HZybEWpdFe167xvyw2tcTh4HyM+hKZnku2l1cLHYZjTzYtVqAlzwgL4q8Hw5j3Up
5N1hLbdTgx9qMBLZjk5KoN9qi9ghYERA/VaKyYYTGNMLYOW+fbooufHzjW+EtqyH
SyaKVP+h7Ccjg07YKfIfmI0QNVa7bDf2foA3WZscH20bGswfaAXzIx96cjRzg8C8
DHYT/q6oZVLQ6bDVIM/REGrShqWMGkzog9TonJ9+q5UU2SyDTpQN6cj9BGf9eq98
llm6Br6UHLPPFu0bDlw+jrB7Gx2HNkfgG7bIVFygcOmgzTqu4jX7M5lBAl7gRzDo
Z3Lk0VDu9MKImx2G5OdxzV0nO0K1XzlnpdhMBmGqeVB9XlWb1hFypRZGowfGqe5P
lDooSZpo6Ipdmr9zQOCg0KB9k+BQgwaR2PxoiPyj3YrqURkKlF8ZpP6bElPFIFl0
KEXtD+M7f4caktIvii4JPUiCu53fXxAvAqSsJEIrTY1fmWOo+fWjzFwnzHhZhQLs
aM9ZEb+v7A9a5u8Bw2v9LpxZ67Ag2NO2wBFKZI8oaagpCzhOavtT9i/CzoM0yKtV
XeWBb8EydYMZn2e0T+dQa/RUpJP1K0npE58oJrBD28nenXYmTSO4NeL2hdklhN0U
r/3+XNzhUUg+a6nDGxvAzhm73pxlSh0hbGeKx0EPGD0K/9edqdepCaUQEfxVs2II
C0wRtxHnCra+ZuBQQG3z2wJqmSHKcocFxiay0C534u0+nhfr5+aYyt6Uc+Ax5OjP
KDqY8+sH9wcO1C7iTzICxg68miXZlaN/h0AemMydj2aOpgiyp8gNf235TSKO2/dx
Cpc9KOTXFQzwLH6ao6KsTGw6bhk/IS3056M9CiuYxbxPkGTG+qxwbE2gq+Kzk9eU
pwE1/xR2eqGC9Zl+MPne8cmLyZ0GJBEnCWvMtucx1lGMguLYfbjrUN8119G4yge8
6cnI8UnVaABBPWFL0OydPpgwszKRBV1WX1/4Qa0oQ5UW+SPh8UmLFiE5SpGxcybu
w739Pr0//IGN0Crdv9si1D+d0Cyk18LdJuWH5LU1AhiVhSBHBhRBtVw2F7ta3Qro
iJ2f7n+J/LqO2AgTewFTzaxP0n99LFnwVXRP7B2e9fgpCqt195V9LrqMyMFETsFu
H0R/ktvo06iq2zOtJ9jjQZ+UfEv3ZWfZuzXJhcBLbcdf/p/d3gKbXdmAQVxIvS8Z
MsOJDX/UtKDsbEeWc3Uk+2W2WxXX3aWwXm0OvgErmDL2anCCzsPRSOy+XrbvT7n6
8bzVuVNbH+zPUPnDbsErh8/Lwt4u05qEqdymeEOpSPLnP+wgholQOOJHjRMNQn6k
NO79KJ5LRc/jHnX+YXD7wuxxU/r/h9vc5IOwKvjoLTrK4MMRrAzHqC1yYFMbR10G
2g0ywH4iLYHUqOWEWH/lhCdP+tdjvo8PuE/ePafempRE9t0Cb25S67HzkUiRAqsa
Hnx2Quu+eOnAxOKSqSuCC1FK7q6sk3IgukjOpMrdNW1yWJo3qv6MraD0p6Ruyclx
l2cnvXCci8QghZyyInsAG1ehrCiqnb+JccRntNayFK7VgVM6+tm3NxVZZQHZkxqh
ui5bh2vhGlDYRhsKPaf5Vih8KotD8CH5B03YAUzvBu0AbvPUerSqh3gUM6gfzp5t
hIsNZxqJidNnhC/jAZ3peY1b9oG2eT9Sr6SR3SAxLzFxIAVGKbnp6Rv9y6C/F5ck
V1oPloih9+NG0jyD1G+4FlGK3VLXv2QMbVTyOx36Ccu3u5vGBXrQLYBlNu6kNRs8
M3oI3zOqWBKA6eoHFNLkZ8TuQGZwteexKbLrRiTyhF1xY2U0HziyMFO/x9tiZvAd
GPNKlGdQnmDq7HAawbxYKXdDyrMV24s0+1XvZRywEoAIM/I26r6c9BEXpLQZdHZS
6GTOS7sXV87CZkHIsWIcRd94uwrhyq9855VWyZs/gGnDyitPsnHUZbuYu0rJuoRp
Ps5pI90DkpwZhP/KgvOrIhS664Ao86J+TTJziXYgo0J4zH9khdGcd4u1vytWjg/7
TiAxJXlWwNrbrVFtDjrPiBWpbEiyoGiTaGgtNQkrmYMTLXQAdDcgzfL+GPIQJW2S
VsxonZmSmyLROyixvIeXuB0QukP7hsqVhqBv7xLgDUbwt2PE5xKz/Xqi3sTTasnM
kgISz6ZwUBGWnuLwV4TbVVj1uNtLkxgI+gFnG6YXXdCV6wV+R258dF5K6jtRUIz8
OqIj7AplZUjmwmvSn6CMhxd2nNAiUf9jf7vC8dxfE0v5AzJH2GOHqSARbITD65uA
S9ABA6M820T7OOqKE107echf5gwKW5aeJjmlwuMzUFYbUv4yLON32tHJTikS3p1E
fLMdrA/ylBKolGROpj794Pfs8+UoWmieFf4KMonBhL7Gd5MoA60Q7avVeorzzfy4
Q/EDQg5UVcbD4aupcf2Xl5ZCXZ7XdL2IOvxcD3h6vVhO17Om3r+XuUGUZHOAHCIr
IGgAEWPO+TDH4xmYfx5ULsHxO3pYpxW8W54yfBtJ3sm2mQFv07Ib+NOngssbaHlN
0d/VXAji1c7tI0C0pakifKHF+Hka6uWnYDqePwMDwZBJtWjlucjOB6TYqggEQZPv
/64PM2Ru4tHg9nlnTF9dYyyhZUMXoIEyfjLBeGAgAJ278/aCzpwDJDo0jes7nCKk
PxRR3+JCaocvGNbe3k02u1nPOM9+ycHudhldB0NMgGS4qQ4+IOJkc5wJguA15CJw
8UjB0SZX2TL4lJwDcJ7bxK4ams6vBZq6w/ff+jbzGS5cXIpvuJjDPm4Uk0oyZxHr
xr+67ur82XUZJDUDWkEcc6uDVgTt1eYVcamqaj769scR+2Y8W2GdlOtMaIpUC1rV
H+I0LP2HQUZB0AJlkKDgbrAxnCvUtzUTlRoZlvPQw1S1SVouMNJmt8gMTUKni/K7
tT6f2AlP20DecqZ6Wv9Qu12VmbR/cSG96/L5TamrLjckXWyFNwPVHIvzZLQgvqIn
3NdQm1HwItfo5DNn1g6OoqqG8c/hwyKj6lEtqRRvEZb6tXQCYvdXp7y9tnVs5Dsn
GCsfJ9QbxejS+UNY/Tn8E3v+fmJ5UyLqKuJj6TJNi9F38b49x4RnAGR8x3+Er1FM
mrzgetFFa8U0zXQ+UlTC70cMiVH0dMJXorYkkibTTGidNvhG7iz6MzoOzDzqt53K
psEgDmqZEO4FmEJjdgAnbfCi7N5GLtkkW1nyuXDOOem1pe620bwTSN5ORVpzDfQ1
ISZN+zhleAREP+4tQtwGUhLNTrdmMeFIw0xyFoc27fjwHnnAMrqCPXxkkLg0uGOy
NAJCrLsO8VEykGDeegzb+mszQkTdO4wKz9xIwuFs1rXTQhYUlSuQYE16XJhkGLvo
xlL6XEtdV7OMdehm1qeHeTuwoTVNe6wyyJeu9lWOVr2SvnW8bQjtUlaQvZ5dgz8r
9LrzdsvxbCxuFokDpS7uVolLVNgzVVKXlUdcXi7HlCg9dGMYe5YzrfGXtowmUXeY
r2GfM5fGAutW0Rmm4flx+j+k0RwzWtajWYUVLXPBBrBZsdmyZEm/sGtT5PHoPFCi
B1Ag5BcHfpXnom/hfFtrdCkdUedUEMGX1ZMfpEXvzVqSrCs09NKM44mkVeCMr5yY
R1ezBU5YCgO52iJ07ueeQI1lUdage1iAEgqhoq2hmqZvEClqmG3q41TTTI+KaCq/
Z09up04To/YN37uZVZ9gsgiK2xg1YhLsRqMKxN2kUaLoW2AvDFM5qvgITr1Pu/0w
Y+MI3bO0xxnYAqtU3xz6dVAkW6YYeopeUVRQ10KniKybyh+bznCH9LOBO4x3PMWz
O5QXhkQ2eCT0ovCCZvjYHUzbFQkJxNpusMDw2pAU0sAV023JJMLGaVejT4T9ciEV
BQA+zY9wYLwvmk21ffHMIDrAyO2sMxrS2iV/ortynr4IH+Ba12cPHh1z/PnpoQ3J
lq6eADTWvjbTwTtAoGFjdDHkqXSRFLoxzDTj+vlMwVZcv1gWZXKhMHiFxdwlxCX6
HEeP9bUV1TOW5fsMOnNoeCpSrXygr/UjSegm+81ZYI5eBtjJscd4Ll43r6Vr83vD
DHVhJ8t2T1KZDTQRsKm1M+4Gs6Ms60d0/J4V8Cm1BY/gdMNStKL2cg2ot2mu+gJD
vmPGIT7lPLaw84rmfq3CXWIqe+26aCBaAbCgxxsQZhAaQyC9i79gg8tu+IYXMypc
KysX+3kV+1K/0z+rf/7F32WtXh2TvcXFHXmrAFKifxwiAq7gg3iR8/Pl6pxmmOTc
xwC4cllOtADgWRVc9/wpuSIX+MFRVfNZHyHnwIb2iu1NaLMvqoKMRf5J0PWALgVC
HYbcfXR8SGZ7UldrD/AslJAvSZh8BRnoDcPAGjuIEF34gjIP6k/T7dHVHQY36d1U
tX+mHGD4jGoeuAcVK/5wzHz9xKAPndaruYLy0+Wp2Jx9hgUlyr5wHCV/7TBwFE2c
4GHeL+vmTEO6cXtUdjy235nlAhjrWL2ggRlVz2r3i5g8ZajFr/sdGqG6oHbZoXOi
9Z4KzRZ1JMQGdDMX6uvMWRr+77w9m31VRIHy2tZay/KiIaiPNL7j7i/4prqDImQ6
e6hQ7FlxcQsRCePIkrjlQXpJzyS6RzKe42+uU7+V4Kfjh+XXdVH99s6r5demK0Fb
xxxL2mi4KwWn9kutHB/cQf69OwM515efMhp4bIJ77bzw53Y9mDjgFw75kqyMLEIM
x5MmqwdP5LqTzhmTXOmJDBmZ3EvzTa5PiCidS8kRuqi+O91PaqbAqxJFfzNuxBiP
XxkETRmsf+hFnCnQc2n5AqUk5Ubo6bEifbG2tA39HRhtSzcm+pvIu4DcmM0YwMCY
qK/qndy2PWBgG6dIGDLO0mtY1YGNszb+u1GrMlK2n5sH4OFT5GfCaJEtM3YAOgpj
gFNkmFpXfJeW0acpowwf5W9yibHQqTW8xWMQlgliTtFLdy0xvj+Qh5sZN9bQsCWo
brD7hsJBUaON3pmzg5vSbcL2NT2Wy8dulHgXBoooVm+CD3HGdHYT0605FpyiOtfp
DH5E++cA6vmtaRsPu2xw7iZgcbjE8M0ykaP+0y8vJjjslN6ZuG4vQp4pIggzaK2f
0VYjYn61sPs7oeckRhdrWpCoOIAtntMQuSZsf3hackhHFU6/j4CyFrYLBMomMFPT
4wbhAfWrAd5GJ+GADZIl7OffRsDmAZG7fV5pgcqZ/iXVZd1Vy5qeDjTzL/W1mef9
G1bzNaBHgjV4lmXgthGn9qlLrQi39pRBQwlYmyl3c+b5go/OndwcGiurlHVTn0PL
LvPAq98vxyz3FTDpEJ3FTNl6hNjX8dqpthU7fm1S6l4yMRrxiuivEMI7u5B6U/b/
RH6E8fNuVILt2P2BcGw8BmkrqItKYjg1ICvnxsMU3B8hZcU1Rjj5mFVdUgKDMbhn
+jxcwOJtQzbrrCfdVuD4HAEofVQUrI8ogfSZJ6sXXCoRXREewwUKB3avdXjhhZBX
M/G3ujVVTojAwnOS+P8mo0NFFtEv4XmDrjwK8noZdU0PjP04gzzgbsE6lp3mmN40
0p7y8hzMZdHQgtoAdDUjBgZ9WBofSxBYTIS+PUSeWWOpoZ9dUNRgsSQRxW1D9OeR
GZzM2bMWq0hlV1Qqlob3XXXitEOY1WUkzN74KYL+Tm7LqudsGxvBoneOz5SCuhLG
sfAABBXArh05J7wNhvEs6Dc9VGgK0qksFoeEgS8NDH8vjIGhllJ6UACZFQy/uMpf
GzRY8cH/PLYFL4SKgtWEYmTUbNvD8si96JYfY5lg+HP/yWgTWQhQkaFKiXlFm+N1
ig4GrvJEZvyiZtJStNtu0FXD3CoRVjwjTQuG0wtMaeVfRYtVDOtU4Gb8/YvA5AlF
rkLo5WHXFWQ3lpRWvQxy5NtP40OM06P6fENvtpQkOaTMjEDvefrPeT4bql+WQZFx
jfRYzb9ysX/QSLdiq2CKUduo5oXCiBAhRP0vw8fkRWxFYiAQJEObJpgyEGsSoYWg
CTkmcydBMxE8OVRq79spca31jq4LSeqGouZe7XE0Da6lSjfHicEt02LVbJWN8iHu
7Eq3qOjGM2/buGjpkqMUSgAidtR0dQG8PrtNJ4IhZRd/R6wXk8w70usV5gPfYt8L
qkpIEXFoE5TlWdhT3oM9q0vbF87b6LRFVRDEhPSneu9+/9uKeBp9ZtetWXajz9vU
jQWUgWmv1rylN2v0H5sTizS36VcY2o3QkIHRIeCHKlckOhzqfneguhqbJyA2GqD7
3zHlMLQzqg8uJVxz6Pm/QPEDDMVBaLCGzpFNs7PeQdbO5ybrU8nD0VX8Oqwzo837
gj2OissGv+oe0m/SCDySDYvBm9Zwhidla43HyEOWqcVWEX+VZhmt1ekekFiuOSbe
3An73Nz5VM8clJYX3dVGA6bw0o1dQzCfj0S5vJuBtSArIhtxNIpD0EXN9nVOIx9p
VQXN5XyGKdvXPoGViASf7hHTiyTrqokmbfbw38slMTahNs+dXhE7oALM77b/VyEL
PoV0smNvw1FWR3Vz4PxwAfwKDRVHhQ1FF9Mn42iq7TB7GigFqQm3mWJuR6GoJ96M
LRQxTXbBjWTlupldp48K9z0APSztxw9vZqnO/x1D68ffve6BXkDXHF3+Mk7q+nSg
r1GcAJNK+/gxAjpfK10Cl+O0veCdzP7fp5LOPla7lJhc6a9YORRBztb+nhCU/30L
ObGZ7fvLgAVkUUGqBuCSEXBr/OfRt/UkbaxEsCAb0I5UIbu5KLMiHi33D6nfhxG+
kKYw6T+rLjxnneA1Z9SyHVlYYIQ1p76nW0Zcj7K7wqtuRldDqjABQEG1SqfNVmL0
6mGE+FGsBxVI8FRiE8jFRLpD7HWyQHS8oZucWoREULtc7IbFUI2AAAGMUP0EE8PM
aOND3MO1Hg3poPyFhrQ3eXybucbP9ruya1ZQeyinplL5jxBwfNdQ297HSFVQRTjy
PoWz8Pbsq8xCnC+qwMrgv/jhEWnE7bULbLfB4gnsCzwTagvKf7myYUXxviOPkbH1
4dHNQcN8+YABH1jWvhDZ8UMktJ5xkdevb8xdL+kOzuwQWphTZYalPCE3eX0hyfOb
C4SYy51Pt0BX29PEgpHrq2pmFAmMvbTSwVKl2Y89nkb5Zqvmam5fEyH5FOPc4gJR
svCz012SPY6LItGOIIFd/wmWNYbX+lxUSvAEdG90zGi6QldS/Y1SfitOeoIOhjUf
z6xZlgJiuNtZ5/TbGyuoFkXrXvlF2AK/LRJozun8GAnWJolBpa3cf4Eek1dPPrMa
3EfYk+6scbOS4A0Ot4m2zIkk7BZm1J7KmCZXQQuEmfZQvK39MOAEzcW2NQJRibuN
DBp70sWdoMZKqt5TBYUGkwyicaQc/CA10XQTjOZIdcml3bErKruc9tYUezW3X1vu
KYewi2bJQ+NDFVThcxn5aDULaMOZVdWYun4ezptgBba4IVxw5S++atAAg+dZueNm
9vgpJkwyRpo4oM+UefkuXo+nvnHAg7QTufjbB895LHZq/CMgR8bog6lIfG9GEGI6
6j1bpstBIFaP8OE5PKdYSQFjSahZCtu3Ve6igNIhNbvFset1BWESDzzQYOQABdR9
wj4p3D9re8PcFBWEgsy2c/PARyRXSQ8oTK3p96nvy5reH8NsKlve6ku6yE22Z/EL
qcfh6r3RQ1MKy34+ylAfGxJ+570Gb7i+ttpcs94v8+WjcmB/iiXoR1somN9SOQZP
C+ZXLE0xBAs/JlePMevRkG9t/ei2GjEZiXmoCH0ObBf/gSQ7zd7QjWhhbv29SbfY
6T8Mmd82bW0ChrRpjiJhS0tX+Slg1YLjOyUft46tNTd1csg8HfJ4BZw5OOfB0Gyt
L9UuYPlIrmiTftVCf9p6NSziWO6+T6s9/UB8Yz+fMEsP5aszPk8Fe+Xc6zFQ/HF7
X4jgXyTsqsfjzjnIUtCChecm23eEstpn++hWGCfZlHNWCTRzwOCUEKngRQLqzWt5
zvsx4vF826wZBEZkS5cM620rsEtPigCSN07wf131IacjcoGFyFviS4PKcwqaDgex
Mo8r4O4b6n6SmZK3XXljYYEpeDvb8PzcgEY7TpknmdSwK61mawALzlBCLMps7cF5
kfhNREjKCy5oNdWyY32RTvOZ+KjOq80CdFdZVt+YBSp2g6RH3QJKLnV6E8PMlYvQ
pRFbag5z6ZM5PuSGkdOKK9p84PNqAY4uwtrV5XiGc2UV/Oz78B1vmDVV6Ao4b/Cj
OXeqjW0FHm0sQFcdJFxvxZblVyv7GunfNLQzU0o7qlq84A8zDf9Z52zf1aAvVlLH
Fr/fBapQlANoTEoAA20c8JTL44uNTHjTs+3LZx3GzTiaDjuD89272I2wNl9QHsQC
hvTPoPmjcvCegpJYr2BdXsPvn1O/HwAV9Br/xvzdBAKFkBbBlD4rbaoczNtPxSt6
OyhrilaqkQNzPOBzLuxInnlrrYX3oNhz9WYuLFL7U5ctTq58ZUg9LfFFQ2eI1tCl
00xzwwXxj+7ntZ0uGI7NTFJf2dwSqawvITiuEacF3oHhF9PjcLQk1Nc1dg5FnnD9
oPe4Ec6Jq96bNSMlAlavk2XsCurhaisSswNdKQeuY5w3oikqOaWk5ri+O6Kg+JAp
F+fzKVTff9oyUmpWK+SxJoUfTqBlf5NznoBtLaB5Rpn0uekNdQJM7TOzP1mfcwm2
KkIQ8hxhS/vt0j0e2YxHe03tnzWT4IryErYdHj8ZdAQzt2ujybgSOtNggYoP5VW6
NhayJMam0LyxevF/cTCdYbC0WzDyQ3vm/Ytz0d1HYPJU1fJ0yehNsY5OiELzBpMc
2BwaSp2MKYJT0AjV0rm/AUj/7JrTbyl8sMoslRqLeJw/X9UQgnKRXN+HiMg3uaIy
wUwS8+uAMVOWT7YGzG1FIYLQqhIasq4DjqNy2O9fb6d7GEFtyj01uz2fORokerfH
9qzuir5IfjKAZfYx+B3fiI8+WMG6sVctT+6aXhQ0SXAWMVN8+LU8GYPjF76JQSYv
K04lYlGawrIfTJnLtDEi1fwxVPoGR/tStVfbgZhKTClyzcLLKQqLrcf+Wp6FSVSs
lKrdp1x9WrnrVgBsn5I2mLo+Hp3cPP7D/onMfhWWgprDOXQWqrURJPY+pCkD4rI4
+wQmEhgTZresZZnNoU7MW42nwKqcGygTF9j1OG8O9NnOQ6WiVYvFJOiRzO8TCzjf
ted/rI+LtrlFKMxn+BXpvYDq5/iYJt/HmX0UPofbFPx/vnN5aOtj5cYYd40/dwuP
MvuFk+PjG/9uaVdhq3+CDKJLX6nqKFOddxYj9Ldd08pn4tOvbXW+NhUq50e58gXk
tZF2TE6mlurfSvZx4O1Bi08NcJEHhR/9y7x20Ya9F1sMXJRDzDXIQZLFsjDRnFz/
srcz0SG+8nghzWUcBYk+6iP8CMnUicQ4Lgimue2/SXS/oFRdQOliL7EznTuZ/T0E
pcotspyAMEbJKYGInDYHQpDR49ilDiySro1Rs1DjnYxZDg2VYQGu46qBT/4E4RIV
DP92byWjfdI8H7XhgWYSUPAK23LRR3m71XA4cD/nh8xzaNYNeCnQCbiM30Acv2Wg
n7xDLUQMmDQ/a0cPsnAgabsjBNRsqNi1/4THfGWz7KfQbfiCofgRT+JvBTbLGCRy
3+J65ozQUQ+/Ea3lmQiWDfFMe8uTc7kMrjKbDy+eKa7DJSTXPxO6Ch1lJJGzwgOp
0uRg/+pzUiEA1dnuca/Rt6NnqsEuDt7AK93/634i/f+tX7cSXYoROSfp26rkn30t
SR7INkldBnMEFwrbYvZyS1hQlkjc+oso3GCpuEVXF5sz/leHoxlJiWdf9AL2u7Uw
7cKpF0zrVz80kDCzwf9TGh1dvExxaG4KoI8HzJh01wPBzUVt2uTtpvAslNdRvRUb
YR8virxKc8oPeg+g+DPPfRrpuEdwwp+4aeZkozXYq8VgPxIKgzio8Di25U98KWIB
wp2K4tU6slIwEerGHueXY0fg2a72CAA1SavlMhBPSAFV7/7+Sz14yFwWKNlZFd8L
ROa+YfCSlFjOMSOojx/gO5RFDJjXDKMcz5LxX5/Oy5tN2t8JscczPpZ113IE43O/
grBUlWSXNs/qJGXrowAqhtE3S0Jx/EqaYLQOU0WtTKGkdHGQBSWbRxjni4yNGhYd
StyRkeRwHu6T/ePziSJ2ufEyLO9+Pkmom2zYC9eB+B81RHqFzImtDPBUxFFo+oTr
yYBZnJlXEdpduQa1eJjBVeldjobn5NB7gxwZLfJIaEd4w0B012vuygCHn6zYcARK
UQz65FT/So8h+tyGZ8JpUEziW+b81FZkjynN9WdomCLCdMK4CzaMDHdXXm6A07qm
86ST33XTx6jc36YLroPo1bpFIVcQ/lCSJ6322iOnPxkZdmBsa9ISjW4Keeumo9IS
ZMJjXMCBCdtsfyJWlIYA4jIIWpQ3KpcI9PT+l6L2YN+OVysqeUhMuWPccWk+EarN
EO2Z4uRHNIOMyKmvs5udRTvtRDsA9yQN1TrVkghMXt11/KPLXy0poJxYLgQ3ZuT+
PrhhtF71sM36W1uTzhaoRhYn12reWqneFDc/guYJmFly984YjbceZBKXfWw0iIos
zbGtsyiXY6FC/oQbuZF7KWXW42BPV+oXTcAUoaFn1n06qzGOfaGJATWRdEd4pKAo
aV5GEHpKDH6lSHH1w039Dfxz57bZRTyyqptiCsY8Gu1lGNOMbe+rzh8u3uBtelKe
i5QhQ8rlETdJH6kn2WlViRq9B9+Jx1aK5t4j+5vwaFPNl0V11LdBYKyyIm0X+hSi
NjfgZGoaEJLC5lxJAXZyZCzJWQzb3j9TRsK7iaruhlFWKtRNnjAdlPQ1o6jyrN3j
kCPiffJ+XbkG3qDTQMPF93+zJdXESAFAvsE7wZs7mpLnBCVU3Awve/kK0Y4Ohkl5
dGTxQUbgMjnAnyL0RXmpyAhkUvSRXpu1nuF7CxJEhpeTMFTzv9C+Aa5jN9ry4coR
em/roM97U/6tPNfw+uHXuY/MVqOad22hXGsQ9swpetl03+WIFf7gbeiUPyht7hS1
EigUrBijAm453PSwapvOjAchp2eOTD5rDY5xguJUt0bzumTKHxKBzZc0mJNUqUb5
PSHltc8vEvx6bnMTLGGy+HAUDtr6DNDr9FrOslKnt7mZa7V4F2LrPhL73U60+TRg
ipWopXOZc8AWSscw2t705yveKvTrRPQL2eDew/hsz+2bVeBhB6+eoopC3KZoHdrz
YlcOhwUl7CZJRX/CR1mCsqFICE1xB+gE0Tj+ZOKtSSnQgSEcYgZPs7Ir/jCof3fS
OJ/Y+JIjg7JHiOI49aX57vVQidOxY2gwtunTwZzHpL863g+uQDED1V24nFOHuy6e
+RJYFm9bXoAbrVWlXFPgCf0ih7bzheyvd5MQwJbBoVUs/4UVUSKxXijGrOX1/80Z
nPP5OeeVPgUUc1Zgj5Ge8XgxiUhKfmtNqtRNl/vSHSFhOq6TjeFCaYTyOwDMzrK1
VTOOvm9YVbUVkXFgj46thQSthsKoDCnGslZBTuxI5CyarDDZ5XRuR4R7xrwqNlx2
4cKg7IlI1qPK+15chiNvXGfj+0W3XQgJsG60t4iGyWPZ+sow90ZWNRpjXnLlwvbR
2YyHX8vqSInkjUWIdH0oEtOVapcaz/uXp7f6+t7obHRJafCymYuV+JAPPxQVDi1T
INasEWvroSFRqZNvhfTrMxHEaZ2KuS+ezWSERds+58LR86vLp48ICItFrKyb2Xc/
uyO1GtJxVyB9uUHiIv5C8I8LTZdDtwjKBaLVTojDwOIu5NC8wg0/qwht3m1+2N3o
gAZdrIgQ4+mc2CkC/Cb5ag1Veja3rkz+SgHOPvb62PIIY5S0crY3SBDaxdzRIw5r
gzDmreNS3TV7Cu/x4UdJTtM0jjpS7tTLsHgEp+ZGL0IlDdwS+qujDk+rh+l0/Qn5
i04w0PRNAcIAmSeyX0XPCtfNS1qF/fTum/HiPNzs3QuqBPuDJ5UB7h4xJQ9DMJxK
bncwjC07qNUACXT+pxuqX5Yw+NHpEyoI1qHVgzbrJMHKr0M8oMIjdZ+XUWuhoU6X
yQXf7X+EEbKsndmanVKILy089HKNUcJiyIMiF+u02n9wu0byyleEe8UN9G/FAtjT
laTFV9UTagit7R2uO+0otqsFp6h0yja8JqnwNz4STsJ/eaGyTcXVbXeW6Keyst+h
u2DlOxzLcYSn9gYCHdSRA6/tZgOeQhPI26OQmcwx2iv1o++U9ZVdySKRpKoAa6Ba
1Zp7QaT9hP+mHC/LgHsnfxnQl8NtwgmZuKBUWtWWcsuO1XO6kyQWEl7OQFo7MB6E
ybatvH4Bl/DTVpJhOrwvLWWPqHnFn8Xas/lBDko4jTyHDDraPrwrhWBvp8UG3Vth
0yUupdB5zpVbM/8u2tRTEuedHWR/RN5otUD5S7hA91fgW+vXbJv1r33nLC9kmxfu
ZxmCIVk1MDAVOPZ7R2tZRR7Hddn9A0ICHwo6E0uO4fE8vs84Wm0FyAujChhocVk0
kcCdzKmC6tChatif7TJE+SrgqI3tPck1I1RoWuZgSGWV+FCFhJgVB2JMW/PtaCjx
o0RX4EiSEjontSN3MnBycGgnRoYnAuD0xnXP9TnOEtL/Q8HWqRXHEpF8cqqYmRUb
fBjmTfjurp6eWsjwLHsvl8ngne+W7lpDf5V0+tANZkwRH/KQGtffcxYctPg5LkmS
fIXH9+gpw3miq5QYmhyiP1C43QYwMdkd7TyjLUD4IrGxP5BzubXXFuYrzbTgqZy4
/1Amr7KhAOnzcybSjsaPBzevMXKQHOgZmbJjdrOUStwKxpepejZWdqib0nxVF9KL
ipeFcFF1n8/+c6B8C9LiyRx3MahRR8rTraLI4YaBY9kiaerLYkm+dmaJnDebQl+H
OZypsHr4LxXhBH5s1rbKAYo/buvZyTzDt3aZIaJnECTyk/PiLNmdvKdjC+/YCBBr
KynmOP4x9cB5xTAiN5l+aMhjwUsJwKYYyW3K1nUf3nTkL0vHYGx8SQprNyq5Yxwz
icO83IOPpVaCN+BdbJXrTteFdiemSv/Tb0MyKFqhhs6Wk2DlAYWNPUHQ77ICYgbK
/lMsPQVG3ZQRgizC5umLe0Oae90jiOP7Fz0z0nT1OGIIzrFQuLwaskXWN9dgI3Om
c8O9Uvc/72122s2t7qfLEShNW+Cghnnfj3XFWiVHIjZ5sel2dKJCQpIj3R1KWXuI
IbumljdrsNoLOHkxQYm6ZDQs328hV9YmyivflxV1loQG8T7KmMQQVOtPZXtXeYcK
eMlFwKLCxHqhI9ml+Er5PD29DbMISG6jMnRIa2JryMfyDzQNPGUnhUseeBcChuGG
Jcj2Tohn1mbGraxfINM2Pq9sowbBnyoqycVzs1nfoFeQ+x2GWDqbHMV54KWN9clF
XN6jIivoz5JnS5XGfr5nZnYy3+fHvssY3h39SozC76+l+Za6NcVVppjudon01Pe1
zhhnglVTc1FhXJvcb9t1Eyfyo/JsqvlumI0tCU4nIAgHxCHoL0NaDp9uZYLA5oyq
CFjDc6wzadCNZKYDBLXCl9/OY6enCwO+eKy8U6gpUbdroX4X4D9HviSSmudsM1/x
3HmS4B+fMmoJaFOWnsp7S1pmQv1VQUMjbIxvjRvu8+CY0zfBE5ufZfUqdGgLU9pF
hYbe2i/cqgokC6J7UAieD2B0/PKzh66Cx2iYtoMfvVdZUDInNnHRndAKFZL4bKsa
limfTPnuifLwqEH/QZZiU/03idnkw5KRXNr0S5ncuW12ofz9Iy8GlPLupP5QVs5M
AfgXny1a+CKYPIOPT6d5dm3MfpC/U8PCd45E98CwF9J+nrprmGnaDM44t+RqdSH+
uQqKJ9mERPeh+EF4ynsORB+Y4MqAfrJbtRaz3C7EsUs9s1ZpKnrgcyxGSTHauwbe
4hZQp+iW2WX6UZJ25ZHq80tcHRRbRAIrEeWlycjvmd3Za7f+LbrIXgOCGhYUR6Xr
Cwzt7KrrQarkKZetEjX/1oOOJX27h8r+09U0KaNQrqqmMQ6fGa5+2x3lTUUiJoNh
VEd4TWWrCv4KpdmLJ+VETYFP8KeOvmH2sBq8SaQP1v+JyT2vsXAQs3dskYteQcSI
HnxIBTD2mKX8jSZBpta7FeZsZT0kU56pwBnWegP1Ppm6mRn3zlOViHydYWI1Pmb6
IHoXpkQMFdDMyxEvBvHSQUzGNBMXPG9vGiMmmRCAAZ4G05jxYMxS3oBYkgYIlipC
CJYO8l81o7hjEwDeWhRfvdndnuJooKTj1pnB/dNRPMziOJLjZO2N0LAAHBZrckso
uV2KsHcEWTckinc1dqynTKNflYWqlfpDFJ87oxCUFn9K9i3AgsZmo4ZVgjdTS4I+
jH5B5u9ih/GTCK4ZvB5/DZiU1wXLaBN8zcqsFvB86dl0mDYRectHZZG32YmlKltd
Oi/pE0W1cqgFn3L2Vm/FtwV883QrwQkO9Xql7lIsHdqDvYfySLBeRngTbWF/Ex/G
LXKb0bQhhs6B5+SIttvY0TN9BwYpB7xnNbo9VDtUJL3gkfk1I8GEuZswb8wzRbWs
cd7x8Hqc6pYInUZKJzZdKuH1ZwQ3NWyrLlDvF+nMXenJfDYxA4YaUnn6+spVCUP8
FLZYDuS+eN1xVNUbPwWYUSHV9q2MXGVZlZQUhjPbY9kdVtj03aID+2Xc3GDyQQ1b
+os+7Tg93/ZD0JMktvuVk1l/zddr88yxLvykXVf1oqHyXKwBfyKmxvWZv/9qmhCp
1WZlEL8LupTrkFKgovogwaJqefLmYIbfpp3ROJxNqKeXRyXbiao252Rn+je67Yxy
Do4HYNyQTzMv/5oKPLcrvOP0wDk6yB/l3dD2/JgcSMVqSiXR14uV0lQwLGIHZ2cB
IQ+/QE8gTW6w/uwjdvBNuc07sOQFSvjOLBFKZ4n2u+U/pK6/W+BTNZct+XgfG2qq
/d1mcGVreT8s72PZKCUncp+8PAzxVa75z7+RzTOIkqMF4boeCHFNJkn07r17rThl
WluM0zkdXs8KQRISVObg+8V7ViA3gDpp48QA/nXYWDJphUbZbmGaB+eU10UjKZSd
VJmvrsHavavmi4yrtj0/oEe8Yi8/gwecx306BVAp8wQxgCVD6tDwV/JrvOjLmYxi
kPFrLV7n/qjE0FCqJjQ30YsgwVOvAeHGlqrkdKXDvFgChhvsMnPsszmqwwb9ZWv1
FqRn/CdTiaNHAZgNAYRdVWKrbDsgx61j9R6xkVkPLvUBXClyqF+EwO/NAvYO4DTy
TY/VoQldv4YURdWCo8olHf/KUh71a93A8k1/+CVkmPU3SxDSf8MdG0C86WSRpsVG
wigagasjiAx99nEMljF1iGp9FaMpuWaju4G+zmaxyTQz+prmSCr6ICm1xEMuMneF
wNjyFM/QN1k+WxqKdAu9f2lxsCUxb5q0PpZ0unaQUnJKdMTyndITpn9rTG3Vw1T5
gBW3GEao00LLNgrOjfr6Z4wjka8u/Fs3GJDRKDJ9oVRTmIF2R5IqsGkFb2Lkm8wj
SIfhcovIx8Qr2FtTJvNHo6VTMbv3mNr0MbEyUzdl58OqQ7HmHBMRjmmPCKmVTOLR
mVkTO3JXpfu1jrxBnz5ih5GQZHTnARKex2pUUkNp3MTs98mY+RNSsPGlAZz9QBKm
NcUJHkLJoqTQMeUDzaj50mL4uFNBB/v2OmVNlEpmN89VxmnqaJjZ79mOXFJgrc3w
C126FLzrtOW5ZujTxiPO7JbVX6X3FWFe/5Cl7/LFCFwNTcMuVJiCRZqir/7CtvzX
sXoNhafmsxT3ETQPxyrTuuMBGxde9F9qXzZUQJ2xPxdZIkk1c+8668pF//8zz0Rf
9snQMElCo/yqhIhkqWrJ8NFAOmfO6a76bLrkQfsTkLBYUhS5t35qHPWMHTRLuCh0
1mMMMIto9VzITpsp1FC+LPVYD3DeXlnLFhebpXBTN59NV0fnPmQ/zUmp9CuLK30x
ZmzP+3+iIj0WloPsXBCWNIWUK0zbh6p1qIyab4/gEN5C7nN6ah+7PnfJ7oNlRPf5
kUsq5WY8K986XKJR4RwPB7nj1UC7TZTVXRKY3CK5iEmfmYRpmVUTRaJT00ngrY/a
rCyf7aaTwAiJ7ndsjO8096r/ypBXXktPFoyBF53Bm9Ar4WV1ViwzbpXOF3UbWQz5
y7OuPjvX/bi5v52sEz1+pCmBLjMU/UoJCoDJljrdjRdpvQr8ZkDdU/1jhfq+guAT
oFkmhEc91qfqM2TliR/O62I3M2i3unQtu3YaUkNtQOuegxUQZuY9QE+YnysFdZ1c
/0vo2VzrlttxxoaRCLmWuj3L+YyeNCANtOdVUGEtTNdG0Gdt7tRyZuB79he6Qngn
vdBrGJm1tJIaIrr20scj3usJ0lRxi/mDVGbkt6+k5Hjs4sFf96Toe9EJ/d6R0+T4
aE7rFWuQ3jxTVWvVz47zMGIFV9lHRxNCkDvK6rQT9uUFen5K68pikV3Tuzga/MPS
wON+vWiDpVkRC2S/4GqMZk7Fn3T9DYk0s+Di6tVV0dZn5E9HOCbG+6PRu3f14FFf
lS4RxmFMetPx45pjQO+jM3dCvnqNEIilZZiP+6yNHR6CSjjbuMpWbFuf7Jr51i2h
Y6FMfH/FnM5+kWsycBKzv1deJC+iauPoHhIoTBmV8gv1x3o+qqh1ll2UBHjdXxrT
IjXEN2vN98KbinsksroP6416DqIps1A9OoVYqSN6bxu0KdvvVBMgSX6qIwy4jD9C
l3hFzoxSHaQD+/vCJBoG8+KKAHkbZfrQR1PO+w3tJZs+wg0RQprcFZM5OjJHmpQi
9ktYRA+7l9qeT2gyFjYWCtLAIcx56B/j3orUF0s7PRMBehqsr4IRXb6o8NaJpM7D
CT2n1K9mmZGJDdQA17juR/GK7H3MSFAQzUAIGwU10Ii5ToSiie/fqvtVJNvgK83C
DuBrksPOlhcll9xYAfd4cnpBedoDaTA1aGuI5f+MN3GqIy5UIcfUU5J9/KFTFbcu
MxFsSH+q+dCzSyvpE97v5wyEejOVnQBsuo4H8FRI+4Y8zN4dfma/7CXo5Uc60M++
BglKRYy3CALVTGMG/SgfjULwCaUH/31ApX0xmWuvX6t0Yw4Gp/CxPBdKOMNZegZL
NCeyCpMSVT/p/FkxUNolXLfuOotv7GT2J24LmUZTt+5QAkPMd+vnXKapmY4OLpOU
s4dlwJyH+jTrhXs3vw7ELLvspuN8R1WtS7vcBufKcI5HbwcPgN2e0tEDYlCnpkAf
KKTYo9++7aCi89jh7DDlqMPV9Zf9krR6tbWtUA61cKCi+QyJiWWukQh9s7l5Ouuz
egIHjPG6tkNPUuV11+jxzMyJ9BHH67bTXbmKZWVS0pgsm7JbBMNVVGc1Jrq2IaY6
Z3pyMfuQkpxbpaCsG6EJ0/l4JqJXdBbjxGjDtU3prco0/e9vN6Oi8cZzlebBCOhj
ke2TG5CcC+oTamZI6NzqUPDtULaWBxi5rY4I8JUI8bLTmMU+/qOsON+DYWWsijKG
rWZasg1u8qPPEzMmL41xfV2k3+ZZNDwT9tomt6ET1lq8O3bPioBiEfxIqatjvvUc
ZkUranYK5ElJG2/GgtjBcxdQ+gv48J8Xi7E6KFlIZ5l3hSRDYdP6/nkeeSDutRyx
Nn2uNAWNoTuxa4YzX5kvNbHGJXptw9Xx9kaBV77jeKvbSptU+oB3SFFriP2/F/Rk
tV5Cl1z2cbyTGE+mNusYrTXw5Auh2mbND/qvgXVnH4pJ/YjzaK+8EpfGTq+Kv7+t
I9Yhjw0vo7hRhh8ZOG3stasaReqLHTmTiAwxb9RQ35mTFTWMgv9najwpkPerqnvX
gk5JBuIzknnQukJveSxOzti8Gt/TnQjwNSpPSHycdl465MnpQQM1wbhbGJHKzhJO
R7rdgp51wwUs/qBecbRYl/VhCP4vamMvT9aONw17+Y+nltUo8b43hUwYGdwe/hwE
eft7jylmONezEPGikww8mpPBh/X784OQ/6qip6bbQwAoEuG9vRRYKgi6UEzQm9dG
s3VtayATtYhQKj1s3WayCy3ysaYZX9zErkMYgUf0FoujbxZKkavI8HDewC1bZK5I
NJZ7MwX30fkVpNiZXQ8tEq6/zW+cbSOqNc6/gZsxpV3wvTTobsIiD5KKCYNFT3S/
FUVpB3gIsw7HWNITiNFTsEKDm+9f4glPfMytEmT8Y+oN2utpVwrMzSuCI6oza0qS
n54QSJZ1vTHnf3xkI9Nfhr8w6RqN12t1Vg/oBXEN7QW2oTSZVc/JEpnSCMXIgg4m
ttpDpYZOH92cwuMNNjU1eWNbGBfJBgcDGF2FCHNq46J6hJvYHAAAMzDLhbW9D5vS
7tv5wxzf4Mqv5h7KoM56BGcwSDHwvgFWPh4itYbfbxUABLNXLpL1WXBJtQOP54Fn
eigaZ6qQYOyQ1U4Vzv5syPhDKJe/Ue00LuXvIFwywIj65nBCEFd3Kf1KI6SBrDmU
pLZutB31zA4kxz3GqGdQKax9qGuqolKoLOvXTA6W1bCBZzTnJULwNnLawSsfb2bF
U4Qcib6ipfj2ZNIyVHDUZO6IwsBmXqp5AfNVKIPT0cpbMvScYjyfQO1vviaYnBMa
8ogFT8yc+Wng6fnun4ZKg3zVrhGu/pY+DgG4X7s7zPt1EEcWjiMWoM8/kzygUJx1
mi+B6ohMxXiUB9Pkv275Z/Y5+CFD8yzGV+VuByVBQLpr6d/HzIernsxf0LViZUFt
7LVd9yliz/E8lcht2jqvzHMA9dS4fU7lvPMzlkIExAotOKANhVWCXzs8BU2pkmfq
0gWAHb33nRHfNhR+zrikohD9W3oFDD5rmjO48Q2c5DmiL1fBVVZluxlnakCaEcfD
eGiruadArGKEVui1yHU9URPGY7ZFmelgaBBBqlJcv2e6ZnUeezLWCDrk3a8aRr/q
m+o+kWdJmTE+yBS514SNrdr0nCd/oafwJbYwnq2AeJrf8Jjj1rA8yzt40ozHv+3U
md+4B1SK6J95ESHBN5ScfctDPF/4Y/kRNDdWoTgEAwztsBvj32HyMp1r9t9E8vxk
YOBdcS0Ac7jiGR51NLOBVmOJbaqxcuhkY6oFBnHnOhu2O9iGO3xASawqxxiKXzk6
11C6DcTgc/NoMwHhqk5nfRBD6CZ2u1bQU93VjFtMcmCz+LbKmCw00kKq/W7BWsk+
vz3wAxqMthGQByWXvx6ifA1kr2dMkBGpz6fzeLCrT5JHcbWmZIiDZsYrU+tGDsQM
4vH1lfD5zIWLrY8f41ux6dg+zizwulHiahDP1PXMnU6dQ5v+hf/AYqrr9zDO3d/z
/4ydfF+Yl5iM56OpUcGK0fU36qZByIC08Ously5zlZ9rx0UEbXwOrCg+WIrvtk6z
CtXCGOo3bEPddOkMSoBux6pE/JpxezHpmili/qxTmfsb6KVa+tmNIvmxhjwxheXv
U8Jc4zGnejU8RUy56NH9W1qckmPiQUgRFxHVqOLXx8Ek7Dfoed87FrXFHjVi3ruR
wQLVKt8nm89EQ/PjAxeavFeZu23UeU53iBuN3tqdgfsbyo/rojF5QjNMfNVKnnB9
V8ybwWRW3EFJ8RZ5ah87FpBUtf/SDgS6wU2dfmwdc7Jc+DiONQE4VnJ+B5KZ/rQR
qxyN0V4F8bEGZ4LD/fq/D/RdQk+ER54hnKSr0/COD7kqlik/4/+XlXtCOGm1mE55
gSvUx3kuhYiKHF1iUBlw0wVu9SlZXgqIMbLtNIzTwR1KM88BZIlaSRFqBCvBTuEa
GQbHXt3PCZ9io0shMnmFy2qX6OvJCBD13xle9+vzhX3Jmq5DvWPVYupKuy243YPR
nNGeQMPcCP8+q3Fw0jwLznx1Bww0ftknBYZtZJ6A/tmHS8WKyi50khPTjQRehOh2
2E5W2ZxK3UQgVUXwYFEdJjVy+a0mXew72awj4rhjbEogzDUJFE2Dqf3CtEQZ0Efk
vEu0Uhe02/mBrlcmYtiWCz7N2FdTa2E9pUSjNKQSHWLmMjZLuxvd9mY34PNaAGkZ
W4ppL7PEdD+CJs3Ufbpg+VxwmPS1f2fWz2+eu58ey1J6Q+MaY+G4t+B2VaGzMPr5
gzVrIof8Wg1HJRaS3qpJOH93fcWMSv3kVWnL05PV3+lmk0OpVThLutxWedkiaUuF
WkgxJsgzyxUl4w1QkKsxOICBM6Kb1z51T8KlJnTp1ACGfykrGPKaZUYqiw0zpzA/
XsGSZVqyFlSGavwI/rsD0CYNUqGhUdyywf5CgrTYlRhnAXDw6sk4nWd/hRxhI5w5
3N6b6ymm8zNlGu1XZ1Wm5Ca7sFDIVR11VeWsAnxR0DuUWDxnZRGc0rdVz7zolpCi
vm/ZZE610avqE5DQAxiVhaN4pMOyNzpxHkfd4qWQ87iy84J8PqE8Tg2j51xvpyZR
LGqPmOeCKwrZof2mlJ1xeTQsj5yLnPa30A64MuCmz1+gUWrw/yCBIMWld00qG49v
5p5TwWt7KEwvj8q2sf7EQNF0A4YwwxRfdzEgH8JYEZDde25Akz9oM7RJiBSMW2RE
urgcPYTWHuWz6pU+BCJ+51tCpws740QjOHDW+LncwT/Fd9dlF3MmziIjcdG0ks7D
mthHI9oCRZrqnAyusFSCiYG2hdkx9Mx8ZRN49uGVjHpMo9y6L4lhUcXt7LXr66as
EZus4NmX5c5FgrOUo0u1RV/Gse5z0PvpvrPfWK9H1UNztxW7bGgOCT6jETkB2vpa
3fw2aTWvqPXHsUfxUTYqlWWuV7K0RvOrBDMi6F3z7jV6xKh2EjwcBq8jns5tNmUq
JEYPfcmR2203YVZTcXZ180DF5I11wiZB6mDhBnPsKa3jIFJtjhqzoAVQ2v5ocgvD
lOF04jXfA/S0K8GZa76Y3jKlXtaY/Fc/YYV9WKfbaPRWeh9K+27WatBSDhBbwp8c
Mvrptc6gVVDwJ+B307qTRtH/D5Q1dRDkSRvvZ/EiXQUdXNvoAmR2z1xW3gyV96FC
1J2xLh2NdqY4fWsT18nTHHr/JboHN+JrrgsfaXohcQZ2FA8k6gR07tAO/1bmqEsu
BeILWeS7eHvsJ6Q4t2v8BXGE6i0CxoybdHoXs4ErXI5v7lwzqCGD0pgpIxhWy3nL
qPp09DAWupQ8HpDbm8B4v3R/gX9TLGXpsa8PYW02Wom0fUS17av2soru5OIYm0xF
xIdD0w2eQQ0icRMYxbh5EQ7KkqhmrQkI39Ym0g3DwGAeggHCTTMB8NX6RMNwznyH
KUq3RNWU9/cc1C0YjkCdqlZ3RCnCxjOSUEGJGnKvT3Rf7LqgNgwkB3Iz9RAtqhxj
MRH7RuqNF9SuBz2PfHaoCUzPqUdi15s713Hp3wZ96j9QFjJqQW7qdJ6ZdUCZNxpS
euNIKTXzrDL9Wdxw56YRf0EGpm1qZJkDDlwZwRGx12BVHOkV4AnNpMSUXmcv5pLm
O+79QoRrgEtMCabIoUTxm6NpHngw1FU0a5fA1GXBPw6LloE08BbCmsqMWhRW+1v6
7NnL4b1hXHqPc8Ts9lOuN8FlR06olp1usfShHS66olycYjHg8NUzNYa+WoCQIk1m
dNoR2Kx3FTevB7vnNBVZ5Qet2xhzo0XFnU6Y2iziwRBQZCaP0ERrZ+vb1ASaHpcs
CuGm28gB5xwMXZ98qV/RktWMIEDtiDKIlvfesc8olh2dFQLRSVH8xe0ag+kX4JlJ
34rrcY/NwtzS+u9g9HrDvQpx10yI9c4m2i0cmDU5AVPnO5Y10gUukCJCwoYV+90k
qP6vC7ATgILcwC01vhvPLI05y5IlpAqA61BwputQF3guGOc/xuJG72uIqH/ryojP
PxkCgKH3gi4rpVArE3BDsNtDiXkIOIZIU7t1liCXzSkrlAQ/fpxs6tscvOV3AXLa
4iNOuDJZw2/S7sTvtx6eQdtzmaHRGbhyPFmQuZ56rejLvpFXBnv3gQ+GO0YM3Hvl
9aK22IkTf2fZymgbvKNkbKADKM/VjHc5a1oKArSwfNGy3ElYQysH7e0d75o7d2Io
AIsEgiE3C5vOGoeCtVVqcxliAoBRD2IIzmr8XMNyC66Fjj+Tj+yHob0+M0Yxr4Cr
8GfTWfWZquF/Q7Zh7DglFk0GYjQ9JOmU1fPUXWE9itvnoFrI4IwCrA0nyQdRDM6w
1DqfQE0tk/0pbTUo8VSUA0zEhs0QWKnMa/KNMaHzaWz++H97XUjMQE3qfgaA9t8F
T3bvtmKx1u148sRiKvomMOA2FUNw/Wu7NsQRYxBZqmKYe9IOJfuFm6NoNI/mIvmV
UXr/PXEK0GlSNkh9eCiW/47Yx6Stut+uqR8JTmOkoVVsk8Db4C77B31f/yJR21+S
7TLqB7gDFBEr/0TOETIpymD3XPrM7TnWroQCXLygGTOciNsD/3GJaHRKVkAviYQO
jgJf6O+l2mN7oFuKPpwmxUyNE4kODc8evk1uklVSgRPi1AUSiwMtdJwnoiOEE0mD
WYfWFmN5aeft7lGsWrOUD4V+xzCkXm53Wt6z8j/FwQfWOjLXFtOdEC3JWQPCaoZs
Wp3a2XrfyFBZosLQIeHU9cEAZ+cAki3NuuHDuFB6KvEUQtxnmWaqfSxfY+KuB+3a
vQXIMhP03LnSegJjyl2iwq8qIj3N+yN4lNsjFbGc2lAKHI0zXIHWRGk/f7vqqQ2P
PRdYPLIV15N3ZnMOTtiw/E0Lk4jMUi0ywZHx9Lr8kZKbcaB39y0N3L/9+r9LwrcB
zbKlS9dIlxwG0IcCedlmAtp9f6DTTSxBBP7lXHy5lZz7Z8FBjA4sx7anTY6Jrc6C
K5tsHPlkEngj+fFV1Mgwj3WQguPchsfI2p9EVFYQvP7EQVOXVjommtt1WbyKTVg4
06WQkhHfd9Q89fa6Gn332Pa3OTfdVE+GVb3nEw23UnkpwVOyU7hyguMot+UiKczA
k7jz28lNftLLgcCckvpiZCDg/E2rKLdGf+QBBT1oIiw6ouhPFMUtFgYwY/MbIhT0
/IM9PIaPUl0pe20xh6i3BVuCi2I79myv6VN6d97Ek0EAPxN8vqlss1DHI2Fnking
V8CHG0HyCRYVsbhot8gcsxmcR+S7SuhStTsXTN5uJ0VnDeO4JxbfZWtVDPBCRU4I
owuTTTuHxPyBAeIit7OqISh6WhSKoNS2bFE5i5Vl8SgE9GSRBksRDpE50cyAJR/h
sN2sh3faIGV0mP4qhUnDAzDq2O7DZwhsi6vhiVzjceaYPunNBoQodQHFCQLKT9mW
REdfYrj4ZvXKeIRoJZRx2RkQnO5EQackOms4b500OZOF3MBnvCy0X77eXOgjcf2n
pVn4u5/NzhldwqL4LZhAyYG8kGDIOMrHsO+wKLcet5qtE+Grg8nKop5eHzYnU/j2
B3MyrCPneQ6WgpvwfLcsDfXR4FOUaEzYfbmVU+gzJukfH0dmi2Yh+9GuTYbMhzAv
USi+FoM+hkuW8Jglp8zBgV/hJotavaV94/4D2A7MqwZ+AcJ7kzRgr0iwd+BD0hCP
oJ9tyIIc5fhifDSxJDywDK4i/+NdtU7vr13EewfazhAjTvoJcmxXavtQN+NVeGqe
h8X1BEBAU+YinQx7vBA6VuCuJvWeGGswdkdMpRZoGWPJl2hLaYsJ5obaflvYcTh1
U419fGBtmmUS8V+JoRn+VdL3GvnxbLiWPXIt86M1k2Uytberd40gkaXM2sLcjjFl
DwKZ0h1MigNYNBGbN0X4N7ps2I1EeBZJtOwaxes86AHDRLbVj7RJnOkzK8QcijFf
zYz2VS3e2+HJpP9EdKbRqEG0jb2YWOuniBeNNvkJIJropqFW44Rf8mfn/IDL52nF
vU+OC0xz8vQ1QZUXt4fzDzB7T87kuLcEWC/DmZUKJFBuPp8++JSKbg3in6IiW1Mu
7vHk/gHXCc9nzx7eIUNi4T2sB9hD/4wavDK14Zu5Np6DG4yp41rggWrnACT+gjSV
reOir6sraPUEKTrDw1oUFEGIrEYdQnorsHVJoPCIWxwhP/rPFIIp4Gm4SwWu2Zp9
yJlok6sUz91NF/XbnzptXdc1S8yuIaWrAfX/XJGu2dLI6ssenrUKO5DnYAOWWWwv
BuTWfzh4rbvCNVYK+mN4i/FXwvPDn0Nq0R++lduCU6jH2sh0mHiAa6FtV/IMksA+
SU0l8ZttewfMYOa06EnDEMYKN4mjyDmt3rbEHHvDBWBtUyklGrleuVwD9w6ybEQm
gHUaBB7l4wp1G7qWKlk4kpaAQtWk96tDtRdyNeUldUnSnVNaKsPEqU8rQiQN8dgj
usClnIlknLEo0g8X+9l8aZRxcqIlF/MioklfMvgyuIaJ0s7EkT1KPgvcMA8i/skH
KT6dWZVzymrFRlam0pLbeD+Fnd5ISPCMDYYk07h/TmX0768h1AaZ9hgAhAIcPxfK
wgaWIqHp6+Sm19T9NCD8tSD7oF9nVcqqrWv3V8l8oW0frCHjk3Ud5CYviifizsLn
HMF2Et56juVvDyxOEQCliRv1iXKo0GwidyItTqyJ/Vt+aSPNiovuBQKA2WYyPEfF
tGvzrJE7Tyc/PBvV2brOZf/DHYB2beuV2NEa3LZiSq5aQJ1RxA1FKACPnJJlKFjd
eQApjJEimogqnwHqitJHHjeq2Jko0eX5lm/mD6cuGtQtgwcgd1mKKfEI8iJXYCQi
bcNeX72R4JVLEjtp52XNJi56dQ02v6UYf2zhN4pXNY7ziYdeKWtjebisy/Y6N4B9
EymIR07e+K2stTTMkyZ4T47aPifhSeEidWVJII7ePaLTMIgXbJ9EowN/PcT0vcMf
77LfwyBSK/nN3lHoujjZjFOjFyd4r4X0ilOlz12+bIeCzXjWaybjt+erBs5R8lhu
X1T5FP/bARbFI67NsjrZqZIm/lpbtOWbw1LTKvt8A80ihBOutPIR+mp2NRh9Nybo
DuRUYcn0yzM2dDcWnrPNjlre4MxG77NgMJ+hwcUemxfQIIgfBuwTWb7TVuwDEu5X
TX7XQEPY6WTynUL9sGhytgbKGOCGpSfU+5Ucsveg+EVpQOipL1pEH+MYhN8J8Y79
KiKnrxRW1PAy1x/25Nu0whZZwRhfNRsPtyEVBH3UawWoSTQ+WMj8uFAysFZoG1ju
F2NCb/lqGfin9q2kgF+Iyd2H0mCtco0sGrk1hrhiDKaxca1hOcav7hGN5TDMqzNt
6fCXRObUbQNWwhmeuSsahWojakOD4SgzgxkLy93TTmu3YcpOaL9YjKIWtO2XMT/c
41Vl17peRVqmQFsxaUds0ouqlBgDUXdYzyl+1tiOilzOeV+KQUUz1ip5pGznOuuu
1Q83lqa1kDlo7Ch5yKMhT+FnGinv+elGIov6CthNR13joBt/zpT5P6V447YH1bEK
XaBlXIoanu1GLKdk7BSSK6u5rnC4uObvCMSTKGZGXd8IuA+X5+jonv0v2XRXUyu9
uES4aebR1H4bl3x0y09OYQ==
`pragma protect end_protected
