// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:08:00 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SCtQMquUmZXHWIKP2sRIgCEkIIsS8HbGwQXkaPx617a8mzBKZN0s+HJzl5E/EiLW
9ydTDRCLGh27eZ1v4bz9j5nrRdPuF+r1JQmkH/wNb/9Am7fFH5vsbPezQBkyAD+q
rB+zyTi3fsytQIiXT+h+Jyh1PeZMkXiqqYYFIsZxQsM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48736)
6NHg33PzUKogNblazu6OYTktIGGv/SjM4djZBeJbaxOe55scyPtW7cfLL3Gw3SUU
RyeKNjNrkFeVAhi/99KIpoAHYPhPq1eJL6edDI00lAiihF7qXET85rZKChZQaf94
1G+Yg3wlLvcQ5yD1ZVn5UkQGsxjM3IPCw9hrbG2mNKGbHUIECFQwJbH6feK/A2OH
WBy3LwTst5fMr7CDNkbIvLMv+sn+dnVbXg1TLom7FHAMvGlqN7fGXqr24Vk9z40U
1TQa0hiv0ybzUMsQYlgvt4FEPsS3NqukYi9K0pwP0lt07FQECWGz/f2/MSNhxiq8
UOw+wtc+/2eVHwaGfmicbQDnm96T0xBd+8SSQjxmBqzNiEKgs8629k3hngJyme7p
Ox7nKsokaZuSsVH0EHnkLvRq4ywDW4jQOYaKjSx1ziAiT+4VL3YzyoVhNViJ2tPg
SkjumiNiImL+JN+QLy2wK/nuZ+4Sev9f7fvgRTbpbW4Y8PuflGQbU5FHITlMu6Zh
goKMYE/1R4NWQSmvh7BRFccZ9Q420dXAhHzsoB1RIeNrUMjUa+tvDlhDBteOqDgJ
bjewRXnuZ3yuw1kPwxh0aMZ8m1IPcOwdCvjERNSCL7W2CPJYhcqgxmuDFcprG5Lv
ebe+nO6fER2v0zPgt+EfVx9zxR+ALRwCmI+tYJ2n023r1si0nmOx4SL0euzrRNon
W028+5aafp5gyH5pmFdK+ZhsUohbaYe0wN4FvqVnE72lWu3c5fq9jIvdbI9lfccq
SzK7YjprzilQGluZ2S1XkiSw5yB5HcNlgBSC+OIUR87gr/s9tMdkrWHyFgm8gLEB
qteU/SLbo/kLUnnBq2ZXJeWN0CDw16VIT8h6guFHAf6hg6Da830aywvpgEsYMv81
ByBf2PZRM9M1RIImUafF8guRbAnLXWDqxJMgpknjAeZ8jMKnKM8kMxDo63F070Kx
nMI/ZdO0RVgE0lyiNaABIgjmXD9uu3Io1DPxQY/ElmN+ZmlESj42VFHcMRwRWqn5
DMp8yr1N5oBIVbLVQXwp1Rv9Xw4JwpAs4zx6hINFnlJ96C6VsRkKG4fOocZX29Vj
9n3+mSJarR9c4nE3kI3RaBD6VJPw4Nt7nGZQk6uJ0Sd84uPi9zPXYbRDw9Xk2RLp
G5K9kPVxzYVnpEqWrngGKFkEnFxRLsGWw0QpQm1n0udmkcznzKAQJk6IG6GWrV/9
L4hv1gSQleexKyHqoQ88jXBDBbhK9NPOjrA+lR440aMdceMcYojplCyz9KfnBty6
UaA4Q5GJISDzer9pKWAPUp5XVXfYI05TgW+xqhGWTNWGeFE2lLusYe7kjYKI4fHQ
Sg7DJ6kNmXuLwaAXiweEEwlSpLdFz/PH0WkLf9BTG/wGDPmkYt/UR871sdW5OwbZ
cxAZT1aXND0SeG9HyN1G2igHcLOXm+rR54mndrHHNnZxfkhklHgZepzwZpIcgpsR
VHg8rvH7NzIvEPFmSnTIG03hkr0YDfRsUX7PkN9GQdkBR+vlLmXjmyUI93NLERHV
p3JstJV7VPOv7UhFy7c8OeZa8tL+03PxhYNfUeH2LcJwzoQp2+VeqwakdXtkpXV2
DZT5HEKIiomHBqcC9T4b0HG5Z+0PY7llY6H7Lqtqe8P1bMxa4bDEdbuhDPOOIA+C
1SXd8ZrKB2KOdcr9mEwSWcXkPY483mcxS3RErDan8oteqn7pVmxvcBnMp35WOv2z
BkFUVM7u78qhG2Inu/vTYPxCan8rg99z3ed+k1U9xFYWge5ssp1CXCORfR1VohTm
/77Q76Q1hHU+b5oBsjvWxTxNnihCnpWku+Twc82C349vJcSLBL2cf0Zu8I2pGnZP
4nABfRYp1zlvvQtrV9bX1G88FbnfSm1WBMTeneCCf1FNjSac2rCVjrUrBMSVbzok
lFZhsGkONQS8iChmjc2RmCrkcA5Lt+exMAVuOwMqJPDEetnq/ojFs/OQC282ZBaU
0SZJZZ5zdop4kU01P9k7hs50EKMcLNbFCO8ExM70Y45ArmWMurnpOBgGVLtiSFwq
Nsq5Gp55+LW/bnGlF6ht1eOV4pj6zdwcQcDxl/qp3PeUPd95kZ+GXOYNZd4kjEkP
aijqH0MRP0Ey5O+kV1D/WJNmmSj1LMiLnisZKeq+gZXkFMguIlADpHiXkco+x2jN
v1OgKuhAKF8nbGLJmkGqlcRJUG2tNL31T7IQi0zmCDXQrV+5lsETPhvC/4DU9P8G
PkWrdWJjUkIYxT5q+L/PoOIHqOn+u/d29JZUmelvvv0EzBsoGIPumcU1I6WmVydM
bg1hPV2duG1gBGLs5oKN2+/2sQ2bKM5tiD0uwDQoyanb/vrT9vhS76ZSPkn14owA
pqxQsuZ4aYIkhgdFbQpixD7rIHsgqPzeybU5E1yKm0cmYPqjUIP/N4d/Gisv5Ycv
9jRVhkxnTTzVNXBjCRd+8cPcLd9pMcxu5qBkhObljPq0PISz3DOk/nGJS7wLHhyY
BkUJ0W6SfqIxVcENBzg2D7etIWD062qme9ENwAkzaL41tiR6sBnkC9nxNGJys5pd
SF3Zi2RdpVFoueDEMemn1wv+Slw2QTypyvPbaQEjaQPHs2UgJCdWpW0bcaASxr9o
3oS1Zw9Wegcn5sVSrVGxUr5rdYnv9Iculmjv5ZNhAiP1avzOhw4Xs6lrMCTP82NQ
F1lKtP2XuXk+oUROgjLt74uIyzgIk9jEM6daN0qcgxxPHOnPViekABVk3ubJvkAA
UuuLfOvn8W0vt5S4af7nqaGeeCUaUrzQdhZTW3M6bWAaO0h8Cq9Z78lj6kvTnQ2N
LVlSRgOeF31GeQOn4E9FUPG/yLfiJOjursREa7YHmrUV7HjMbJG8F0aa8SWijBvZ
E854UiD+l6SpwhmEZFtssRlWy2LPuejKBlGeQSrVQnhy3tEiH9tIigboWePHesWZ
BRo43T1GI04nwrgZ+v2kdxYciPUoPbIVj7oqZeeFLAReMOfCXVm09/PiGvlRtGf4
xn6l235AlnJTHPda2OyITqJLnxt8WTw+8g8YtGm8IsUzNCJQabbxJwbqUZ7ykHZH
j4mzFKrhToZpSEmizBKlQxMO+GAcLVvSfxYYTb0KRzZZy39Bg/s8mBcFTq957kCT
cVp1bmNf/KJj66d12HR2fGX8vMvUAc7Ke51aNvlaq8cwiVp5eBC+X+LQNC/0R85X
rIVSxC81T9o3tXO0uivaerJXPOP1TdUaYxxnM0VXIL6AneMqVm02/PcmhQRiBsn2
hDnerdpc9Hp4rPhCo931G/a7+l3fot9vjbghxdbIymT5sv017Xa+nVxf7rIveoH8
UQQD2jTSl0SGSru2FSK2SIRe3FVUdNBkBIT7hUYPQ+XNrzYzBlaJywUqbgADcDLu
/lGGXaYU9iwTKVhNqUEOuTikyPaaEiGqzJex3UyP93p5wO4NXGRGgP1Ayv83JtHd
M1H9PM/QxtCzS+tde2sYiQk/me6nyCJVYF+9rx9SaBXdUYuM4znogADfukDNCfHJ
wSa4oKWpwBpmLpEVttEX9PZoW5aBGPW3mLtJZGyr7tZAqE2NecxCoQXCka/MKG6O
DIHzycOSZQW8deX0yg2jZw2a6IS0AwqJM9BavqPz/zi0Jl6P7kEGFES1DYBZCy3N
fACgCDzdMHy1495avDWPMPSEIxaWK3gfz9vRm+9rfmt/f7VhKo8nwLj6e0pRIPcX
C/cYZqFEATwNx52zh3ZXhdIRJZbRp1qe7ifoDdhzin8w/KOS/qC0Y/EvoizwjxzJ
4RuqqKX0ce5H3XoiF84WuKGmGGHoFs+Bdhm0fbTesg/r6k9p9eLS3i5wt4NlJ8sQ
oieW97E+Jpl799xblIl8+Q9i9gobi/Kp2USd9ZwfkN04K4FthA0U6ylbB/M2cXWu
S2CVMiCuHERGcuyCaQARDZ7c5pj16pdEylUb1k8g3OuNlTgZKDZslCyz0e2dcB2g
eQsRzXcKLl5vdvk36pP8mlZxbhJQcDxFiQtoimMNRfMeH7AHv4LqfAj7jIxJbJVb
/Co2f0ZUJYW+ibClRhQpgnkUoI/vi2lC4no7vEo0mJXyQX50O/w6jXhNCb1NXYPY
i2OkSmytmWtOk3j4sPfIXOF4JRg9CKE7aH4eVk/ccMQk2+aoIoy2/y7ZC90VDH/e
Ku3emZptG78bNg1DvwosHaRWR2XeQEqEbV8930G9epRK7dKvZcrZhsOmjenficO3
SFd04UjXQ8IAMwi7yv4tO2owRAMeUFdM/ic0Ku3gU55jWf/ieRPIlBDVL6EBbRpf
nRP+7+UKB8wPoS22n4QQUAqcdCyHtFQY/NxYENIZ/52WmOzExbcwr/wInYSpHIiJ
m6GLN4Uu9ySg9ZCz0C+3xwFQlYy4yaY98W/TCd0bAHrAWIjUPh2jzsM90KwjdgtL
b4fFlXA6h9us/rPX9e+qxRsiulp7WMJG1F6srjGiKx4SnDjpm3UNYJ2vgZrJPiVS
5lu2SUfaShisXUYo0NmuYgQwdK8YgC2XUqMe7hwrVwwQD/DG/VswO0nw8qycxST8
NUPhHqe80jJljvszumh7JnBOY8gKgZISAuk5K0DchaAgXCMhNn1BmHjzR2UdgM1V
kdlgSBU8XP3yzWCJBjJX7pelfaCZsO44+eWLH3hWUPziiAAKE6iIWlkYjvqMoea9
46lZXdWKFTb4gGsPmWGJscSz4Navva4iJ3cJ8JzTdYY3nJgNgs+IuKJNNo1klH5r
poZY/ITsfhnFgg5lvhTbIdrYw8P5+kUds3TgebRNU3fuO3bcwpCwVEYPhND09l2k
EXHIRdBIKO18GE0V26yZn/qwGNF/lq3G5m8ou0YsARFXoVuYUAh1uYFecMf3f0RW
J0m/FKqYNbcW8NCuSUjh4FpLWKtEVj8hmS6/4yESM7vOS/9NhM3gMISmnZh0qbRB
6W3FpB4+fXiMPMqbFJ74aFE25x6CInmVRYyeZ/0KV+OpUXl7NgK5ON9wJKm4KoSg
sZSu1QIIKTgCPSoZlN7oKLYmIYLRa8CGUwjEIb9aJVD/Z8bmi2QcfwOBp2DH414x
r9xxpEFd5luY1RUyFMLQln3Y9nln7s5i7bCRS7YrLHZNb1ifsqUSNHMB7Yukh3Cj
Pqh0suqLVGnGjEDD/6rj1MUl2eZDRB8qCSX4Vek8JTuqr3TcyeNoB7noCwwcvE1l
LJv6QNdShp0+mora5TMMtK7U4tYgVQAY0rvbRh0o1ipbs3I2uqUMJD5mpp2flfbE
I8xdwq3cz05914OCeE5qsuvxHOKfp/HmrJnNRMYDf+cexnoXfy8xKa6bddwG/mKi
wRdLBV7PYWrSgiJ8ISIsdLU3fShK6s3BCbKoNRoXhP/HCIdU+o/E0/HkgPHdBb76
D/tSa624YrQ9qydspui4BVlv8Yte66y2aq4YOpA3BwnpEo4HTFDp+MKTqwvv7khw
E6BGZCBvWvmDERbQuwubbz/fCDUBVbbhvdgwbZMXw9wEZkO9OcSiHbksdLYEMSCJ
XtUIMoG+X1JW//47XbgXGhYJGKnkhoHwqSJ9wFfK5F1wDc5hwEqnTudl63aJwIie
Nc/T+52O3WCDG8FqUtoJEje4siSBfT8L1cfz/dWn+1VY8RtVjRb5GhiYgiV0PANB
tkgpmg4lSjqC0/oNBeXWg7DwpOsMmLt6F1G/WSrJPnILInyuIjGsNsM6USuN3kG/
MwX1zrpADycyhRYu4KPoOu6JagkjN0SWxrbP9WKNM6GlNnCtJM0hRzMdCewttLbr
jfZ8xA8/KaU2InC+/v2L8wc4LkTPxjoDNIb8CWlf1g/HYcQf4kyqf1mBT+iFzLLb
u9rQDa6UJxo2hKiQkZlhMF1xbg7dCAuqyqW9ZtYGDdhX+EgWjoolUnXnR82uH29L
ehus0SdP3pnvH02Fa/hT88AkAa0e8VaWnD0G+Nt5pkGAhC2W42eYHfwW6dkyWg//
Cc3xa4PptaHCxtcDY/FXLcyNL8cBvYpg0Wt4l6wnB/THRoUJGh3086vSV7QCx57B
Jrl0P10up8YxPHp/vmFbchspS266EKHZrmF6irWlIBkVJ/UHAhMQQMaRSKzL2Z/j
+Atkl3A38CV+qiwnkXH1kb8NaMHFG+TQ7bwUZnI/d8A3J3JNNPl5EGKsg2s1CCde
javlvsSleYy377t5Gkx7U+m9q3zlmaeEx1miUNNCZex7F++lkLT5pnsiiP+ogCM5
9TQK1FzXpCp9Y4kLnOKiQZJQm+4Z3JOM5roBiqshxTGMhrQhXI+iPrTG2PBHfK4t
v/69R6myQAgYChF7wN9kXJWFrfNDqroxjKwxR9EbBskezNcT2/QKqHqN4nwuYtQl
BzvilJVLbVDu2VGgxDFSmwmOVledSXVdl3mayp257pwgZQollemar/FbMPh8BEZt
wkrQ3dWFMzBB5zK/qXwjMWanx/pBdpIlSbSN9aJwMFZfFRwg6o+yHdYF32Z9oQ20
cKEN+U09GFzh/LgfhgSaBBD0NudOZiRawE+iLsyTbmzqqUz6iHvIQN1UuXGR4FBg
YH/JQMy/hgengeVgeg601jDB4Gli1Bp+mabzfPs9Ea+UUs9QniRAXo28qhDap3rm
tJVNAuDlHXQyJip/lnLWlQpzvzr8NvkK+eK+zvr4uzhkrCyJswYuRvcE7WabZzrW
7O106XaWnaT4zCSfr0tFtuNnx7nLJXjXG1sAnlK9hgjp2YPrJrKyOPVvgBPn0LQu
tkteoTKuhuRH5XkeMqp1AB/15sbkPxmaw0GX8vZ/CB9j78E267YjIwcG9Wsi6Kh4
7wixLnDtrXeahNJzB7SA110PAy1Bp9KqiCH+Umal1a3ER8uzt2mh8Qu4rGolKBgM
7smANL4WC4wxGhRId4vkg6QxXZb3N/Ch9lKcg7Yi8Q2byaYan9vvlkewkYZwFu73
7YvRkVJApqVf32kIDv8kmPOHjDsxTXPjpkz3W9JLp4GVHU1YavsuLSlIK3htzHbf
X6rzDA7fDQqJG6msVgEaS8T0revBTmbjDZ8EjLHv9zlkhvQqDwuZ/It6L0BtwL6K
U6PPPRkT9+JLDqGIKwqu6qmTgWgS1zIAKNsD0bvgxvHY9nKVTX3twV2n5KTn6TLI
ESj4T0lNZ7GPwWVpzkAOknFE7mZlM4kLoPRlEi8xpLrqrrAEX+wC6040WQf0Dl5G
Hgy9K0eXI33iyGWwRKX1vnHvnaKoINcrstr3bVvjHd3tNZsBZR6vLtVob2PZjl/A
XpQ5ikIgcXVKN7cjq9VS6cllzvg9iLcXM3Ah2lUlS4UncDrqmPlUKNgazzeiAzIR
iFpnRFjxG9YDN59WSzQlUqjdi945t4nij/z/Qydd3xTTQ/+CoBU7nZ1JEPRtxPGN
NkQqnU9yftyn6vj4qwlFZTgimEXlDrnt0zR7p4oBaIGMWocKdYTIwQgUQaCg97XQ
X+dEIm6pFydiE1qmQVIVcat0shAlIlFpXbmU7vfJx20Q/sF/4Bc4iceWUqssjVJ7
T85PeLEsMQ6x5tppdV0am5DDfTnYj3B/SSFEaN7zmx1er7k75XdbVHorWybhRUy3
6ITg8JgbxSy6xXiJeFphkrQTBhPXez0MHjianlY736Rcrj8jISbyPGOBi9BvQbu8
efKmh+kp1qlgTMLm3lT1Nge7MjCGfoCPvrvwVPVgAH2Lv68on0UC3clr1qYYwOFn
2/PIVl7u5Pi5TRajj/luQHvMth3lgtI94+nHjnX8HCr2phDFlWdeKRr1q4ZB0OoO
njSpqc5r4CxLUAIIKxsX6VwtjAPchGmaGgDUjxi3JAuzS4CqX8mZrLTu8kl7TYcz
jAnRmiKllMtFDuCN8rKAwrGz0N3oJ5w3jKQmILA5lqeomCSHyB+cCrQBXuju1lQP
n61JmPk3YAM4iKNpXAtAMZRHehFaFx2AUIB8Exdv2Sf46VDTsg0TkLu6jkEyR5SN
iS+5y5SDyxxho+3WqTpa7capijjPn9Mp1xWs8EyXUhGosuN5EYsZ7lmMyIrKexVt
u9lCWqXd/LLhXkA4Yt775jKfphjDwqyn1oDqOxzg9cZPOOz4AIpuORK85XJkTBLP
2Gg0n79vuEAHWp7FFYf7dgnPjwtPn4Hv4Zv4pfBfsPtbER6pJ/zQ7W00ufKh5z/L
pSwRz1/2ytsyIJdRF4xBji/c9M/4KrBivBd+JHn1E+NcIGZWbWlxxUvEhsn5xlgD
fVxK2NHKkrfn9XZG/Pc4xLKPcdPIG6ZIGTCvOfECdGl+Hr5SeQshUzaLEvo0SDLJ
PhfobEJfCEfAYhA0ejJCuJATeiXYXQiwE0UR2s1CuxxITtMvWiOfZRviPsDOs1zS
f8+Up0SX26S2UZnrsfiVKsicw2ipqc2mOIY0/YxCbOfwAQtatp2zdAjWXKo5LMr7
/FaWllzPX9naCNfEOtKZi2QvW+u05JUIAosQmemHl6N60qdVV0JoP+Jz66RvYxEo
DeNrH/Zxpc24GP3GLOd8qpPSTJX5NZTFpZS8mtr5yfOVjlcJfirU2E1pDE7czpEt
ObPVl8YiZkmCp7veWnftojFR9DnFbcfsURMSWK3s3nMCEJqoVllnKTI8MHiAlPxz
vVjHb6dMNGleL6O+002r8GfXnyS5Hffug5MOtJmF46bNFCVJBOmqh+8Dx3LTcZdr
Ulpkkzwin/SEH4fexJwOS9ofLZaUCLtC8/U/zol1gearPfrgZYeLfpccO85xYoD2
K6E23bUJhr/w8sK12pkiGFGchBeGFFPr/GDxpFyC6WGktBJNi2DMaBKn1B7HOXLw
NQuIQY5Qsq1DP3CnXwFEtsFJTJ86DnNP95S9+D4BdfL4qv258TXeR61WyZUzM1Wa
vX9OjjnUAq40lPwjtEFmW8zOSgnvEBCeAd2tL8L0uI/XH1Q7yJ3o5AEoeGqf7Bih
5ACA3HRtjd0nU4GqJachRmDV20z66bJ9QrowV2JhBmgQpvplZfTFR2juuAIODQ9z
XFevFpIlBvA9fai695A0X7ydDhN6i9N/uhUSoTWqGbre2iKTlXzmcMkF/4xkiuKL
IZPu5wdMzCi1tOmHMlltZxQvr8WNReB5tOWiggUPiO/PfZKaTxQ7ddsN/kpFDYgY
3D0xJVWzK26YedJ0arHKieRAT+NlZom9wUR+qtwhV6WAWwU6Gnsj4I6wQpPb9dK9
nl43L6K9Mzxor5KodbtaGipiIZnggiakGhy5KXmFaRAJgdpbSTrhZlmdmEoobQR/
UHSsLapI+kri+Khs9JH9gw/zfX6zoLbrmxD3rbB+o6shbqhoTJNUJ96ibkPkQ53L
eEYn/0g153kPic/hVqOBRqeb9YPGznnSIIX8sn0AhI8LQTPzavuJEslWSWque5oe
sXpCph+WSHTQ+16rD2wWUJlSuKw3tLc8ntPwLoMt3HfRtYkUyAMvmtHYwJqMgu68
ps4+WA27DqCtlVbEfCITqZnFTE97mY4xEQq4NxPy3Ug9JCFDE8sMcjHIiMMZCn3N
aM5XMfY1odkWwlKZniOzOel4P8u+3+HkZysYy1BBKtCkTtPgu63JYmmcQnCKcg6p
N4HNbg87A5xgvUsi4BUwRGDtx7jRg7ZgKf84ahg1nHFjfdWWahqOoxWuGBtMXvrA
sWoRlL85R8Foslu/8SZfrpLG2EaqmSQTqesSY3Woi45e6KNXJC+WPrQGT4kIsx1V
pbzEtU2mhQjK5jgaxKp6A5NjpXJ/x2lkPI+Zi7QY8YOy1uoMdans32QOAyRj1sPg
LgypXVBaSpYzhw7IJz0tH7COxWt9V07Br1DpAF1nEZJJQOD18AQN2mt2OBDOM07X
M21Q0aVUv3zd+IoeLdY3g3Z7U6EUN94gCCxX0r8Kz5Rn7S++bFy4GFYu5Jf5WAeV
0jf37jlgJB03eKhATv3lbqoPxFIKEMJ1PRQTPO1tLD5rV9NmkrLvJvhptTsHHrV1
Oi2VzA733cI1EPVBUe5GTKDXhmDI0DgvNqlRFg6W+Wryqw/VtoSxnIkJqRI+PC4X
w2LhkYXuaDPTJsCtjys2MWanPKUnonnpChPX1+H4gvEccjP6gKhOz0ZN+oCpKiGQ
iVpb5mjteP3q+BAxWfFTvL6j+2RN+9qR4XWrj1rJYiasjwKtPiiGF4yeOOQuJuVP
+uDUHkFdFlfHlU+1kOgadNQJOxloeT9VVXqMnfJsLi6cDyFhCCjE1ra1dDWojera
V3rPMV62KHWC0qZBi9QHX89vykHHAMc9YFgcFuZuHbWK9dnB2ZbSlxc4O1NPBdcy
IvgNcwlU7UIhAt41gfNOacoXCrFb83kUMbsM7UneCG7jIsZiZAlORyYGRI44UkIC
on17K53UHPzw543oI/v1fjLobgypqgTSvaqCWrq2h3Fr9pNaCF6/KZqKtUduPNML
qCjz4n8o8vX3a4O34iLXg3LWhPP4USso1+BlTrybSpweiiE3kaXRG8yX/QnWmYYK
PvDLKuaAFiy39BOO52TtoXUq8w+xKG+kHG1GKAY3mhzxbL9M3OiV4B75f/gO6PL5
PppIy+eBziIMlFNn3g//WnI2wBtO2iHdLYl07P2ZUGJS+QePV27esbbQDPjEpVZK
VADWMt69O3DI+X4Ndu5x4P0+igp70ggvKCTIi9FPdArslWRQ9rb1C3+opToMGhZu
Fbed/QGxr2Kxk2KAruk7Ob0Akd66zJTBpkwLs4iMfazW1ajNYoOLw1G7gnmtrgjq
JML6H7HD8cUapQiNZWH/PH3UJb5CnOQOYp2Htewh6+sQBv8feuJBa4IXGx1C8fOd
iY+V2skDnkV7UpGmoDpWpaWz6y9pk2mNnFj5QaLlmrNKybHtbEjFRQJmbzVZfUFf
2/Bc6/LNFQrrk+OG2EBIeJ/c3AglGuRkV9hOStKFbWcn5v/xfCgi+AecGO7SrwtT
48L7cuEf/c87TQcD/TjuaeoFbVqM8C99nBrcGvn8XAXZQKRUWF/b5sO1rfFkiUND
EqsIpVopKRnv/O12ug3yKicXiOAvdICMDYx7mcE/Y5VPVHqkEMlRImzJvO2eKS9g
BUzrlJfH9fz+JYwc1jDk+uoUWOtwtSXwB22rstn2KtgmuBVj/pAOkTkxHCT2QycY
/Sfh27xRWo2mFEuys1JkNE6Z0GnKaSAoxHRe/yxjHtWouRRXzWh88yuJ+lhYU1FQ
2Jdxb0UpCRG0mnVURzx8dacDokubuSHfh0UMe3wSLX24V/vil3x2419VcqwcE9/G
whx/SuLOW7TOeQ/T2GS3Vrs7mXIHAdw0Pgh1h9a05g4i6q0aFqGEbb+T8XxyRiKr
/1DGMbpy5QJBkjdHRIW1WFqUwg9AU/YjDddg9wD68CcVMMxMwMNwWDA+qmH5i5Wu
udADRzHy6LYKD/vvirDbUbtqyf1iE5277A1zp5muMiRmDUd7+M/XmjMU4kkb/4No
9/hGU8fw8Q2yG96eRtRKF2bHEU1v60te38LfbXquwhILmKCsizBTPoZF5U9Xhhcw
QfieoXwVrbwA2+Mjna5elHJfDE0EyFZR3YYQ0TxwHTGUzYzMlK7mwhXmgft7ex8j
/9cQx/IYtzmNaWXNa03NS6uyfWVMqAuF0NS8uysWw0boQInmM1nPbPtexYUIlXYh
mvG6PPe8pFt7F40xZEhaCkoeHZn8z9OuLi0szmlvVfZ7EqhkzpxEjmQj5SDTbftW
W/0eyR0ALV6h155QIJCT5BhDVvolZRMtBwxTa0+7IgS3E/ijDPFuZdZ/rdn+IimS
yLIho1oKJWG02XXIrQQwTZm3HnZVN7Ni2nQ638R83bOGrybjF9/Ne8Z4QGNDXauK
9xmYTwSeQZHv7estuawmQaAXwlOX4JNbN4iIsg0b54Qe525NRoS9sCZKBU2MqfLT
OEC5ReFDjJlQPxUFd3qko2XCudlHygB1vdIum5jEjaT+6yZ9Gv/SyK4uUtWGt3RG
3fWK2w4yP64GLO6KRq9XkmYEjl/qbShFQPN+S3FDSoo/jnE9w1qmXlu/6wpeiM2a
AAPDwNGI8oDuBEVobYaOaoPzrkfy4mhtdnZ9ocXiiUnG9RfiUuPBO+qP6AOhjzmS
h04GGOF7laGEpC2wBcoSyYaTwPe/3zCIToxGTp7ziL0J3p1y6ef7BuWSgmvTx98y
zHCjB/t+cYR3mLNq8CISB9Zl8yVvga3EqSy/8EeoYRYSuRwfeAdjU9Tik7A1ZP92
gqk85Y7xMUXEM8enyFwk06m3ajEgXBitSNf+wN7Fee6ub2m/udToNm+q4LSpj3vM
jzkRP2U28JRpJ49EL+0uPc/qwsP5tM0DC1qcNSc95AK7MpU58+ousoE3ZtOiGIQW
M/rGo8d482j00vEO6+Ed8htAOsMB1xOwOva0grZm4IYgGx1SbOLw05YSI7ZiC8RM
TrE9ZjYuHLE5GRx3USw0Cz58Y4uUtFQhClXLArm/HNjMMvJPUxAdFfVYJT465gSj
BHrzMD3u/ucqNo4Z024wdr9F0eRBZ8tKYbj1GkA0p7+rmRd2apCCplPdYilWisxt
Cru8JkUsck0lXJojlwWk24F4RFwPyYCh/a/ZiRm09WutZLh0cOgg1bji/obYGIxj
Wp3aeafeeqmClSflITeCoZkbtDiLDuPa+njgGuPssgbS9EaHg4kZDCDUvgJLowB7
i7uE2SBlaNrL+vnuM3P5Rn50z3XIyTiRFNumQSvFlCggdYh6rskhavDqw0zaXqhg
G3Z1hVKLAj1Gfcca7oz4f+rn37TB2N2ddADtyDbAmG94zviMvhjJHOMUVkS7V9tR
bF4pEJvsE8d7Hid1RqEG/eq065jN/oEf1Rv6cvutWYktnVOwBaYgEg16MwPWSNAu
AQKl2jB+Xe1g2hFNlNjVUmyvQ3rtWkL8xDkhJ+3Uw7XaEUuhpInrdygTpgBNI9nt
rzBDZ8iExqSEMTumGYk8SzAcRRacWoJtkVfjSsitzw83C5ItdQi4LseMqtOamHN6
IW+GZLAsNUvjdWSXlrsFZM0RUTJ1T9lGiAYyO2Ej0zdjmuPJOAy6i4k9U1IVPZ+H
im1Gnob8hHGsFyArrEFccIg8obceynwLYVyPdZcWeTrE15NcRBb+PDFUepg1jDsk
dLWY68ia92uxXFrUqimr1LUaQifdD/s1fjRg60Uowj3pAPIhcF63c3Z1kgDTD7U8
703ls0kjTBMNNm+VchH7GxHvNC0i2D3YeEy+foJFkF6OtQocUkqgMUA3KQxJpA75
w1mCW18cyQ/OSvO0uEbvXHDEMScXg/0YT+RdgQf5f1YfXWWbu9hDMX00GFzEhhm8
A099437UjHDdMybQ92s+SVUuDH25cGGk8rkLnNXGS/kOwj+Wbg5sKhpOMp3n9SmN
2l76MVKTtKPoZxep0OI/rct51hY4rwxZJyGzuhR8lx6nAXUFmQx0p93d/ZZEle3g
zQbbOjtDPiBkpxYomTjQpX2yyROrqVllUGaxEzOOn7TzETErlYgPDMG+zUwzDUvT
XrCZyej84SdDQvq9pFtDf46hvzyRGuHGxQuatH4VoflDjAxSyHxLB9vb321YZLJq
8tSPYfubB61sbqOIj+TzOhW9QTVvLdwNWuIbnEUnG1P6lrHZQ2rBwlYZV0MkC3rx
DBFa1wNQB0Gp1XzRahj8DEEEzMzk2EifUY5Box0HeA3EEYffyq/5q22aMLeYJ2uk
GBonWMTTyDQbyqo3DkHel+AN8NkP8ISaj0SC7MBajklhSDRbWVMIZ+IMqF5yf6rT
4kkN5uPZY57ynWXBgofNWovffYi8qVnpCviz7uKR9BNU9zGJFNOJZQVv2EHfQ6dw
76itrvlZcMBrjsl4uult/O9857NlDYlwlXCO7Z4tXTxphtfXPPQLv4XWN12Uco+y
apk4KxHoDAMQEZ+47cR3lCF8kOF1JZ2URlGUi8dpu2XbfKYwjsd7NjAi4euxPp+x
TUlsqDQj69tc3mysxhyYE0z3T8uQci+BdAs9fL2ysk30IRQ6bH/HmNuKWndD4SRE
Y8e9SaH8z2JqKro2WkMVGFDwrEHmhuoemtaTcmowWd0phouf/aauu5SDYOCroZAj
K0BbKCiTxS1DjBj3DPeagb2ARxOwtRLET6LsvPshzvq3eowEoop8b8irALXnTXj4
Y1vUjyPnAwHQzRPzRYiFYI/b9Xp5oPUgoEscLvqEAg8dWvdRJmTfHrpDWBbVT4lV
HLH2xlFOc0vG1XCHE+pm0IcWhyFuGBqx9c1nPAkDrTBP8q2X59O/jUi2/vc77C9P
nfExdy20ABetZujTPhShzmt8EE63UFHlxPV2hJxEIfbCRm2PE8XEkdnPnoWSNqDQ
GyWeMqe0HXHFRZjbo3QCtbIF9jmL+gr9F0BcFRLeuaEtqGAiTaMM+Sgd/wKNslPN
xPTPGV9PcocNkgZrQF+0CFhpH5mul7W9OvUvEb+vqG/VVgxPYDJBVy38Dv+/rgeE
6z2L2vPXRT9yOrhokhcMmJhuVZI+UmjJxFEpaWRqseyymCJeBKZ8EzQFiq+zE1cX
vAumyqRvXz0ey5oe6XOLwqKnV0Ww4SjzFMDV27+zMUirddAlY2X4bBPCDKZ3TtJB
xU5h8VRrpbhvHjlN2VG42xjyMC2bHs5ylV+ImcEtLNcOsMtF/w7bzW42T6IQC/OQ
hh4bLiTo/kJbF6OFkw8RwzXkIbcZSAsQdARyxPLQtlELmJPmcvqhcVsJu9xSn/TC
HBpTcLMPCDd5vrp8NAyt7Fb+vRJTOaAA5ayA1VE8m61vnJlwZArH+v9ft+ZGAsMB
0jO+uXiK1p35IjqJAid8XaooH8Lb3tpIz2lyuiTHU2AmNFPVzSlMwyQg4GFOTlsj
UDf1z9jwpPTQ3d2gvpLYspOLVZcOljtsoJUEcYsZxnGN/5h+V8gtyxJODkTpuI7J
yLfcSoOSVRWi3RooLrafkBFnhe8y7yfNbgPTGkjZJh/kVqGQOtNrYmbFi4IV/ePt
Tp1nd10lebYiBcQDyFg7wvX3FRHFd4NryB2YUx8b2wXMKZrL6P0Hv7YWWlDoqrlp
8GIzZP6Sd+fUDDfbNxtTYCw0ezWKiiaMp2utWmeBKIuUe0grzO9krO1vx13F6pf0
UCD7PleKVX6DWNJdy8XXoASl5B63VKMzfOz1DozyEmneemV5Ih1X0MkCAWZ4mW2k
09FQSWyH8Y9fBt7EGKVncacRQsx6SssFcZnS/WFNmThVDUFXKCtb80M3riUrIfpg
+ZjXPC/eL4uNkMGYXXq9GUFuYabioWxmjgab3Z8xrROdo0Zy//oRHJ/WS7lWamwq
FI85Nuur2DtBSs1QBqMPPJcbdS5J/dWhWnG/YIuphO8QYPtZf5tbl5faYkMNdOXQ
lO9q0XBAEDDpu+o6GLZ9lvwSzXiHf2crMdM8dx1iQn10IUxHAvoBJHzf6LS9Aj1t
ISm7s6Zm1+vMpTwuw8p0LwXJrZ158BfIvgdQhaeGMEaD1jHMsP/qSnL9/OsKsn9a
rQqYbgLr5+8guV98MZ7sAJg6J8BCVv4ewvIGVweW2AHQQ/X7E1LwxKKNlzz8n1HO
WA9ZpaAYIL3lVoYvWHeiTdkTkQBbjE6ctTyMf5KOjsSwc80YunX2MgBwwrHPHwMw
XpO0XTf4Q7eFpl5TQIsXWjwl34Ye9sOkuYYx8o9MjP8x1yprdAF6uV38XyG5mmFp
VtCEXIZEQhjkdOV5pIMWJ+PNAibjVHkiHo8OoFkS92EWg6GYYpWDgsQtMLhz9FX0
/NTFu/MvQq20cGZXhgnfrm+wHexS7lxQKieJqG753lbeZw12QSUAtO+l9lWf78Qa
pFmLWC+aWItAeDQ7xF6UUJlvTKtzie5J+9kNDIK1pORHIdlByz/lc8bFrtn2XFlq
DuJ9nDf34hkGRDP57cw8yOm+f9UQIhMQRbbR0u7103+n03f+8Mi5daV95qrtbr9J
ktJdB34egZTvJtf4r70hEQNyiS0x2mS2GauQ3xZbVkjLNq094nJkrApi2nSOnW+9
Y9DenSqoRkqALUv6S7b6y50P8wjH12Mv7l/yRxAAPgKmFdACU9MiLN4xRvhEw9vF
nJxFzxlNWPpsBjSxXcq2v8hDMLebU0xCKAGOKYHK47U0PF7WT1V/Jz990MJDf1lI
bNpOQIAXl0p89sD6GfXXzYt0OBHNMLwTtj2QC+n0G7jhoRsnGWiAOQ/81j+cJ3zJ
h9CZ424Y12Q/Id669d8tqiTQen7P99lL7AyXgMB6An3S1jmgnRFY6uWE1wuCHmOt
ZXX4aL2+D2p2zIZURRT0c69tc7rVBTdxtJ5F5E0V3deno2nZP1MfUjG2K769Ycc/
w1WiV/PhtjRb+h2IR4xqp1D2J1VhQIdEbuy2PiYZghareZ3gxMRgr86GuwEWuq/D
l19g6rcEypF6hGaRpyjAjjb6zdmmUBb2SB6pf6gIh/AledxIHeb+6e28aoa5WcGq
s6Cgtzv/LIXEUzK7Rf4G/GsuiofmZZg8q+tRm/mhSoAy7XnKZIfYqMKWYzKem/d5
jpqLtJcAWAPSgQL5vHYCi2qb3+iVmOc+4dgfiYDdyuXcNC27Jm+UYj6I29d1e4Fe
fPVbKVLj7mJqkM6bCnMBsAf4oVl031lk204VlCN803h6MnFfQPYviyfQoiyGf0q8
J+z9QowhNuRkiojLqG0n1vzZmrkuSefS4aRLNP0TfTP0mkzct4NiYuWqjABNV0uu
o6z1oyaipxBnzmIKELS98jihvrgzVnpMxzLM7BH4AQNaj26EB54Agbubpx4aWdTh
/ATKaDE0B81w4nrE51LvkULymZvyLqDJ4EKKEoxU9EFsDaz1XrJRWkzj7ViKnUhf
mSEjsEejQj74VMOdCt511SUfhZTNmboWIaM2jsEl2UBPr/I0RloZ4jbl6Kyi2bn2
FKRtf4OTK/96lDO7xIrSAFRErOF+sxqpWfBVNx5DUmuBEt6bgnb5z0snffugYyNu
KJURFnQ84MQ9QgX8ckU2TZMZOKrbOfrlO/Gal6U82FwXJ7rIpgNAqYPHC/aigzVf
mgJdb6L3n+oOmVgJc80nAZ4+ko8n7C/4zi4BfwfcasO2blAIh4wwxMkF9mTmfTHL
XdAe2L4Vb8hC9LpOW0SzJL8hSL18VuXzmzryn6l1soas2pAqLCH/qV7jPIlr7JcB
XzspfDGHnmpPdGd4IuzEcwiSkG/vLIGmFVsmqDPYtQIc5EHhKHCzY4OVIya/bkRF
o5nV8BC2ypFL4YKvRXQO+TfQPbfzpplzS+VkhWc5h85kAVrGiUQ/PdOqvHsZQgLl
ioKZsDy024mqjI6qJvBa/39iUAYYUNAXGp4uxX/hPQbx5kxoxut6ufI0xo2cUEHy
FdgDmM5eO07cxyhFZwzps7YEuBtoEsfXlHnsSL9pfhYXue19lpSIqOKGFuKtKIEI
l6/6HtufYF9/f1ZphGy7cfN76bNv13RubwnDmVPfJfY3ziokAllNUnqW4cpC3f+U
1TDuzu17Ls5bLWCmr2e7Ww4DtCo57+13bgqI6b1wutWxJJXqK/U/7IlF28xrEKcs
D7BmG3ofG0STODqIlVHoFVeic33/zpFGHbJ4UAM4Qv0yMK/vu/dTpSqZCwrjlGRD
X+UNvQQJx4f04JcRN88Z9WcO0JQEj16WXZNyj0HqVIlWGYETfmpfHgiTeyrYHWN2
t9sMvGSuXRrpKATFe1hhj1qpxDO/xsSs/V4hHdNprQTEsaXEio+xVCzAf0vmPlbz
UywpBcadVrr1FbGWa/sQDCVcOvL3c8bMsiMjPb/g/JgjMxk9j4LRi3uGr275fibR
IS4ohXQ5jsynzusVU9blnI8JAP6p/6g/tH2YOoPQR63/ETCALuRDgR53FVr7Q49x
xzK+Sh50twdayWX9FVBLJ5cAHtwoWpGKZEtEzvOewPlRvBRriyon9RafeAXrDygP
HPh1A/mzgue8GOudjkHdpmmG15jaKrq/EGRIBogWpq0uu8MrT8osK4j/J+Vb+Sex
DvvIuMs0eyI+g77TXYk3o0YRS6+NOlVrNzvWed7ACnunRcy5RmBU3QrT+m2nKCXq
WmrBmxy0IiME3oEhQPzMDCqStcj0t3vQedPVWcNy4mJy03tcfPKPbVOaxksm4zLI
vXHwWOGhIg6kHfZLEDMkOdIqtbROOUNDLYmnan/aj0snSVmYiEIv8bCrm8h3VyoQ
o6bVsz7BvHYh+dSYFwI/ahyy8iSJ6dAUjjaus8w13vKx+rfi2xiWuU654f7DAdjl
sa7wBfTZEDRDAfUabjeuILXAl4F/6ndJNNt5MQnRV29NzQRKDdeODT7y2kRdQn/l
UOOd1L8UKYhbnuwnNOVUxyjQuGCsqYADO61MCBhzOmNdCEUulLPthhQqr4MEBwRM
uh4z/rYGSOXZ6XdI0U4HHhEJ2MpzPrqjCW0YjFpykVlsOCUZLz8atyAbYMP5zvnl
pHTqLlzLI/ADyKRX3+/WKCXvksrHU++fw5cBNJpNTOA3JxkflPzwFBbF/fM/VjjZ
dedeRP96MLFdTsF2Lx5qQCFx2urr567JadVbl/Yr1cidjONwvvV1jvSJXPQLUgQO
L/rkFStz8+cuTDOZs+kvd+VLbYgqXIcuRx05XM0h9W2b7Iy/c5aKO3Ml7xrsNEeU
Jn8PhuqVB2Roklg/Jj431HyCQQoUCXkf9WFSoKV0RSPQ6bxewL2RhSbaQbBYkPWo
i/YTJnJBpQ5BmmND0zcgTcwQE5zLXF9trgtaa5JypjETLCTxXrH12XhSboemkv7C
pSFoOoWyZbUiyH/oVFK3U+V/O6kwXyGOggwvnFCmz0AfBOd05isnOdsFzSm8MYsO
Iq/Bqkt+eX+TVaPsqVKrMTSnL2D4ge86UbTXH3JAUtzYgOAxif9T06p731+fRpnX
YLzpx9NsFxPid/jyNDazLOl0TZ6JLHvobDk4fRSmyhd1x2pX2zot2OolIM+XqWyy
DQhMwJylcTXnds8TAdblkoZBi9fTU3Q7GdJgyqto0MrQQ8fA5HjF05ecCjq2uJYd
KjDk1xk/PmlV3Uqp3/umPA+XlLgZY9V/AGIxa4GwNMbzkXSr8bDRKHx/1wORQPS6
PHWJHJTsnteVSltwqWIdGdFvHrRY38ihRmP/fCFNgZNWsVjBl2Az9vBBEyy3bHQ6
yH8FqPIywVIx5CGrZC3rDUwg5DqSgeX1tHB4CjbiZPjMOv1MJBKGAqnDU88bi4lV
XmR3UJEpV1uYapsd8N5lHRqnRYK+4l3jOsYA7wObz42Afz0lVFvjbDpRlOUgdlwG
/YKTkssBPANd/OTfm8Djiy8AFVcoBkSgBnpcQT07TMgUDKiHvOfke+1/oqZwV9Om
yLCRDb7p83V0cxglhJ+oU2jzKQabIVfB41a/KANftgOHYsvIjnDdKOxGopXyR2Id
BKsay37hYTidW7y/4nobu1FO/4f6/Ko731FfMx2n0V49H8OqEQdqORxlF99SNS0K
BppwDDiU0C2slmCweS88gQNF9bI4mluYYD910S1nC2WekJxKW15OwsmJqO7/U28N
0eludx8jUwhNhTppbPiKwcls41z9F7pUh/0qQiU0N3CSrX16VGwn0SnKQLNw9ses
aKjNA4h9PQJ9OkG5/PZy7bSc/MMo6E3Zw1xzn+AIp0Us7QDeIsdyXjdjgEuMXnEu
aE5MhRhwc9xQY/We/1zC3zECCWBhzUWFe6RBD50/FcVIqEyEFTywuPTQn/0zVGt5
xdQEzREs/FClSmtX9HF/3PuNA7mjnzvAq7OH/T9lYva5cZeN1U4q2ztT3LlJh2jX
b5PKRORZv+aW+Q6VWPwU5NsX6wkanbZL4YuDRMh1pf+fibtWlSTTZbC4x4sO9ObV
P5ec4u2aguoty8C2JZ7Hdhvle8XQ0z7JVgNtPU66iJR+5rqJnK8+cGG7qUxDify5
3Iu0nnVn05+EpLK1KGMbS4pzSuQvVNajp9GlRRRbINl20iQUkzYF0UMUVFOMcr/v
t300Xkb7av3R3cak3zsqvAk1TT31mgLfcccyWQJ78LNlmqu1uCGWTZyE4j9Pvf4B
3H66Hj8yX9aOGHWGbIHSyenMgVfbXgSmx+C7qOfsbIL8bVVnst238Fyh7i9duEhA
3KvbCA3T2sohblqepyLo8fxBAUzOh3zBt0MhwPrIdsm5Jg5SfMC/oUtgLyRnCdpD
cF5Y8OKbgnoJxnBtxTPqhGsF3c5+nPAr2Nvgp+5V2YNkd2HhR2PgrLq/RXDb74JZ
5CFkK8i32JJ2/mSmNFu+jWcv3rdGxu2LQ9hyjw6kkHEI3eUODdylGG7O2E1Dym4U
4tHGEL45ZFbH2/V3PL9PxLxN4XCGzeFwx6hdeFoc7b3keLMf/Aqsp1eDnpAdrSNE
RLqueWLVnFjNyWXbHNcYt4oscBNS/hpVNyXJAWS6unJLvXjbXSEneK8boMg0Nzl3
gRsPAU5oJN8UpFytgW1nicEj4dTIQ5uAArLj4lAmgjcDkM2w017kKahEGq9MpDOB
hqpXjTJvDZt7V2pQdgs06FKu0YTVSbEQ+RpDKT0Dlem6pTZZN5+KhqwjHZkD0sM/
/9UUn0rtNv1/fnbuE+DsbmjrrZbnLsYHLgn6+sstRQCMBsVXFM5cD/sdWv/CObkC
FSVhv/MbVNdEEYca0/MyK88TQ5JABnCOxhotRNLR/XEhLBu6yY/rKgn0l0IlBEWf
6B8jvGlgPJngmTPuzjhOvhUfV9G0YeqxkNRwLaV7e4Yq+L6T3+FzIAB1toWcrNwQ
2jwiX2OOz8Ds/YL+MG1hXQOIWnwOjHbMEF8JNNTfefS2OIyrPEUnhXZ0Sd8ZJoRV
MvSSbw3/HgHXJMBlZ7C8BoQ1FGvdOB8tYPNjyP8pyHnSMhqTwRrMsNvNt/EHniZt
uwJ1tS1i4Dr4FHCRIH2F0qKI8uXuHflCeWPL6SrmjcZ3+eMAXHdjRRHXKpzm/gAB
Uoekgbqcus5+7Cg8+NUjED9/gQgtgUL7EOtzJ8JXkOFhm5Mx/7vUI13FH0/zc1iz
9dpgLDFPvKBmmgRjmVcNdqGJJDVqiuKG3brjSZele3UXJCKkMr3nasC+L1PafZW5
mcvgvQ6ytsnR+73hZ0AFYGJNWmtjwOsrfwoVBkxOfWjRQSFKyPD+6+azcBwVXs+V
wVFG7VUYWAVow5kfIsewLcrUn0/GypB0GeeUcEIDfgxSpHM1c0b6zCSvGdbib92O
1dKTKN9eSALYsmWpdqjQTv7iVBPbhZbZpiTvNG+LR+gKymUuhGXNJDzkoUYABkpG
e76kxfUBPjnEI/j9Ep/YxG3Q914Y7mO2j0Tbu324PE0THto/eIAev/Uc/SMcvNpA
F6F3mlJvUt/fRU74Ij3c9fb/wJ6gjcYHj7T3qPJKllzr6goQhKAkbqGGjKMWmMF4
rse0JMHFBRYuyLbOw+5CD7yPeSwd6ET/OkzuUPj/6sg12e2u38+EmDBlQxxv7DRD
AYdTHC7BnYq6Ytgl3RsCguBXYYkn2gStwNucXuhi36v07mHkqHZIdAk1F8ePU7Cc
xXuchxVvPjaBzht40cl4m7ZE/9yhlWzJPNq+R+khbuUx5XlV7KgZeki2YgWIApCM
4kwuyVf3+1Hrca99mTJArrI96dExkCgzcbr4YACFJx1VQD07Ecb4GfIO3SVonsEW
EZxTFrmLFJZDqr3SdHkUDy3IeEXeTV4k+ZgEmAy52jVQ/0qN5AjncMCPvoOihMHJ
cirWoc/UAPWu9jlRHXpuCkphLDcKhiyQLpiWXGmmySWSQz2nrlgY2+c/Sr+XCvww
rmPtyGEOlusHVKimwTcyV8hbi1W1dCfuMyEGYuTn/OwBxoXFVqnwvslLgNdOArvs
vIfSWmLimUvabyau328BSWfzneNSrlm4GihDvpYcmDqIeDHurPmvcGiLi2wetzZ3
Ro3b1/TAPDlO9jQm/O+ToAXJO5yR4G2Pzkzn/RzA7zpo7uwWmDIABmiLUY0KqffN
cG2KG3bmLRkDhO2dUtdNvo8dhfz/nA4T/M/CrFySxl5TZWJqD+/Jtqs/vlR6wTHS
xCOpjL/0MtS/iIpFh4tervB8ssUlsoLr08STok9qISSJCtqfFsx4JB9ZaRqikmqw
ygdBXnyYwNz0SkQAOudqgfn/yBL/r/RUHY9IFw/4YIRS2jx8PGwccConFQjElEf0
l99PL+RbbhyfvHRvfb064zOkJFZ/2sqcQcG1FyHPITAdLddU7uIXMYqCQ2TY77tJ
pB57kjQwhFan7HylKikNfnTh4mmZtpajWsQQdOJehcccGKRtj0lLcTP03er/GZoH
sFKXPq+PrU6QjTxN1m22JjaZIKgjiOLCDKqO7iAP/Xf5XGeBX7DP9wiyPapA0QEk
kVmNLG/f1wtzNKBVCsjHgxDQtFKKCIRv4RVjZoRrJM6XAFM/K/VQtL3aqIZPbgQV
VXYpHcPJ/CDPrlTxUyBhXW8mWj4pxRZrHyFORXdQl+hhxzX5OMbl93+DI/Vd+1bf
8RnMKUJHO/5uWpiCfN78bdC6buZ5RepLYJE55ZlQZMeztIRN4T+BJ7N0a91VRttT
6CjYi2nPoHx1yg/9kaaBDTNN2qEM5ZJS4h7BQSwGLH3t+NrZXAM7zTiNNiTzkzeD
Xoto9WxmZ5MlmJN53aeJhfJpMussdJyCXo4JBT3CC9bXagj0DimmvqYwUfCL8IbW
7uIAkM0iKoAiowWkFweQV2hnVlNDe5vONyX0F3kx+5nbyymhUKcyzgofHulnggs8
J2lusifvri7VL5fuxo5jaoicgYaWE05cvEpsfSSbpdzi9myadNR7aJ/CZeITj7dL
fnitVdC83scCuGQQl67d5hKDAPjF4W+cGWh044Xxkk7qFiR5XTrodlGOb0X5+mjC
jZMbHhDEGR6Wbdj9Vcc2O1YiJtW+Q8dR3sk9Ej7sEJZ2ZuZSjobiPpdZx2VJig4i
fz1jpnf15eC6cnBVtHAie7kBKeJdObYaxMPNRLrA3YfGvOr08tVwoaTdhCWak1St
pBqxLMTck1BsOh8truQIgjPZG64bQiai9XQlxL3XOuUsDOwQgcAoovwSjt555X0c
C3zF5zjrfFMshH9Cu3gDJZ3H8duuNs4m5eJkw2kVm/MDvbvX+m2hWNE3IGJjFZwa
CTHu4wy2vmIPo5rENlXvbel6XoUVpjZC2PvGF+dVMriMHa3wxHHUdCkMG0vxW56y
mLTatVxl3tVodvB/OjlODtav7g/1jVZwjoMsxi7ZWHeMb6GeTruU++rtr3OYcpgl
/IlGeEsN5b5bFAs6JiSWq3EM2kfBrWkn7MubNcuDz76Yq4rzQaJthmiOkX0nixU9
dzZL1jT+7S1rUQzgENlecpLi9gNbX7sggW3R73h6+6vfeTU8I70+B4b4Xk/78MKy
EQ4sVioFTQw7EFlzYzedgxG/8Aj0/FpsiDzBJvB26xMYeu9N/BZfeQDru+3cSpdi
y/xFPpTANaLd1yhqAcb02n+ik0g7amGxkLmccFpVUajkRv+dC3Nb3N7QrHNlNbIB
hYGckf19E8FS270Qe1PdbIEr9xuUkeIO1k720mVMjDxpS+pG2aUZMrJv0J9SP5DW
vJRkqpsN1wqQ063aDYKQ8oohBIG3sCQ1uqokPqBSLaPboMdhxMOZEDGQ0WdDsk+7
oq/uti86+nVv8hLnup0HHJOriDjHDnnTK4Rwf2dJBbkUnBca9jpOBq31KhgBxZXx
xJ2GAODQJPPVAy2LmnRUF9kcg3ylahBaJmE3qBRDOq8ifvMFpYnAjoR5Jw5NcsnQ
0OA8z8rbvXVjltVTvl86uvnJv1zqF/YSfOzXzauweytSLuQeYRrkz+TV8oAfLAZm
3E39CeefnfFHQBEX+YTzX+ParDnU9ae97IMK1KBMhrFmDC67nuVU07diM+zWklj3
sh7LllpCqEdlkA5yC6GXW2AQj3/niX51UxXk7u+WsXjgEnMR44SIY72BtnLZmOny
guDfTofAGaJd0oZWmLQZRgFQi4r3F7g8hdXbAgbZqEcfnSfMUssdfOoJ42xFhNqH
1NQUoDiBeIm4RrXmLZoenkvcbGOazOr122+3gTqVbJHuy7CM3d9mRDyLnVP4+Eva
sYQ+128VHCHpEQmlgRehK8O4+zcZVXcABNixLlOGrfhqMBPKSglgAXnEygQdgXgD
Qg62F6CIf22xulAIjZh26cT9v8v6jruWEkWpvLzkp8I1JDGpMpANq1GZQbC4HWvp
EKBXv6zdLCG+eWFocQYHt4ZzQ+BgLzakD3CfDG+6ac9SK4fkmeneXRoROgAGE6uD
Hw77Bm/0+8xr4/FbKaILWPEvevPZlG3vsFdfHF9jyfkdBYh3jdz2DXwXlDR59ENy
j05p4Qet/34RLwDuiN8GiugOuQItH765laz2pne8KxJN3G2/o80/rK9iL756ctPE
ju71YmGGjUeQhloufsqVaDlVWn6dEr4zzyqg4I+r7Ye7630R6sLsv3F/2atB33rs
n6X94kfieo+IwP++Tz9G5bBqpXIIUGV8aP0+03MJZlkEZPV++UwO80NIAgiz9XbS
ILry6Mfq6yK+fJ1ixTzv6fwEZ4UUan3uUc/zWvO/xyyOCkus7CW5ij3hDQ5uIb3m
f1rIa1j4W5UQNpY1NVcvjALuithx1nFFBqaM6a4BraefPWdve49v5IvIw2cXjUlR
hr+aGf3RaWyjR38JgKx92nmJRdCeN2vNksV0tlRWqqT1jdUYyJxShXCuY5utuSea
mhbfdf4dZ59Mb8T+GR6CQGuNI5H1vtWNoepGgRU7tzxcZYAC96BykmUiCPWd7sGB
5jg0M8anVqKO3irCDo/8PIKe0C6JDL3vzGbwlsyqK8zaFxz7/TUf5US+73z4yB9D
ZcLpzg7CRcpuCxl78IMnWVcJp+/IlY1rDiAkCVebeCJ6lA5hjrIho0K6Ebe1pBc0
g7QoApDiBVgnMr0Sy/PnU1xsaIIKGCgOM0LsZS6crLaAjtd9uA1w3ES89LO2MawF
FZ4NxhQF0BDJoF4PVkAKFNbsyB5hz1doAcKIdP264C7StPKavQSY7ZzP8s9q1VQ9
VrIrMeZRk9DTypAKqpcUmGCwxVk7yhqcPJrWNTkICzhsavNaxeUiqgwAmXENnM5t
a0pjEmny88k1gAfmII9vghR2e6TPcAD9wPj/7wvyQ45ekVyRdVFoZkRGb/zZ7z+6
mgj03s2i0Dge8j8V8sG7m83sw7Jf/rF16vDgdGmpFl/m50VrBlnC6awptpBU/9y4
ROLdNWRs2cXx6lX3YN6FG87P5XzO6UMibq82uDy3x7XS9hMr5SbZfepnMxE5A4NQ
EX5IUNSFoksyy6MCb1DARr8ljszx/rr0gEbbHtATNSvXSIspHOwdTbkrSAPQ84sw
xtaav9zE4EppeRUJXG7UrJXET7H/FV+7QUjROfA3TVC/sBMGvi9YW8PuJ+s1leO2
y9Zo4gTwtyNv8tmKUZGKuHqybuuS3cZq6Ifvgbjt/Hf4sROckt8xa5oW4fHwy+R2
tnbQTdWQLmvhp3cxNUAqxJRhihQ3/VLR2pE+OSbcbHfUAMpreeFX2pQ7lioogwfZ
RFj+/g+r6WrfJsqzYBtJJ8w9zERBy3oVBMVxQaU5KNoCSRRdLgn0QzxAS3DuIAII
6KmjbWaKwRaJNDmzIT16p51jRKYQBUnp3zNe1o1Vp1gEgqpNDVfEw6MyhSXXUn+6
nxVKyXo7H6woQaXZ0uyz1CQAwqo/VeYnRsoGD7HLFXie8IWSGFGDxQAddx9tuiNz
ykxpG4R/N43Qt3bfbQxNGcHkYYYnwPAcReSS+D9ScPhwFVHZiSnPKsGlaeWWX+b5
x9ZTzNQTJvgLfYfiF12jJF+1+3lYeSAJkaHhUthyVpAB0clOHL77zq8b2qX4YE5q
g8UhqOD9c3GoM2+tY6ccmFGigKdNTMjaAgl+KcWcq5LnG/9gJlNbogSG29+m1Cd3
7+ES5WrQbhXYTQEN5xhpKjPJ0nIwT0vN99qE9jY0+1pwwJb8lZEU1bSyeY/k/feh
64ztRV8u+xpfmdqNTeRiTalZLasLuzpby5RWcNlmgU+V/4jDzbiHRpLAaXByZBI8
d6FjHJzvh4w4BfTJg9kvQmOfIIeJrqMc4AZ4brkpH9DiMMZmyxp/kUyYXSchydVo
Wv01b6vIMD5beWoDVl1XMoyTFlmijv+zjePZIsLuS6C9Ic24guel+Mx7tQMJAmnw
ZJIn2nqiwd50AcZcSM88dKawnGAby0SlVEJPZ4ge/T3+jKlQSGH9UbN3J4lCtXBv
oG6fLUS5hXQS26xKYxnS7+1+W55ich7O/Q7PGInBNLeeivoOdbw6Glu7k8dsxXob
cVXQ5xqyC4K4gatGuboGU8kr0ZaTrUd8zhemO9viEjMI2JjpiN1o24lCA1OdYhef
+lzJJIes2kRb8OykTvsZi6YSFBciTkJHEX+IwnQxSQE5SGM1y7RjiimF8IAmHbkp
kRgSCxmAdiJnDhqQ9lUfTMwCnJjbBt/4f9JukscwfBagwSdUv3G6ghvJQlrHt/yr
TjXv0SETnCGp6oCqcMCRxsvWHCZZvJBUvuCzyx2tFFpRp6nKX6w/fOOXxTlAiX3c
orDWfGLB/tHVhzhmcnSoJ9DK8PRy5PjDQd6iaQUJsevtzLxpmi8qWuREhaD4Zuwf
kGH7z8NzpUV88VlWsvc1bKjWNmEcE40fyxAEHOw6LfH8VEVQk8JMtdBGuAF90WAB
4+LPjz38ybR+KWojs8W51ckyM1q5dMElXI98drclC412JPttyJzPRTyvhvotZe3c
+DpqnTzzS7itUT0E/Rbvds8MIXWk3bKj3y+u3NJxH3oFD2TC/bUxxsvTZbHy4SWC
03UK8gp5XvUTBVjtQmaLJscN/Nii+VnWSUZ13t0T2PiDq2+doitDbpbV6mKsZ+Dl
eHkqU3em/X9kAvdLrr3Hfh6mi/LC80tCiqP7/bkBZzJsMDe/cRyeHIQMV+OEvg/w
Fpr5+hnpbLA52ojRlJlNMfw1HyIxdSWuxh5MFH55Kb6C24zkmbcid6NyNsW9ETTy
1e5SHlNihxPp0JUc+GMQxSv3LLtYX0O1CohWYDR3FsRZL/DBBEZPrzTyQEiclfFf
bWXFLafx+86ZTx84QaqbNhwifOo0EIbIXeQgrucngdqybEDLvrH+ssKl57uPyBtw
8FJ6btkjbjEOeFePD+GqcVUsNZor1wBw2uJeG4Q5ZAEVRI6mfkDeSbeLfZAKVwue
FNZu04Zq2a5CXEDfa0zWcS7I8ejUh388G/++KdBvBbbowod11fbkqxjEvIclk6fx
Rv7PI7tYPydBW97qlBRgazpHi0Sd3Z8qXP+u5Yq6rEYgS96W6XpLqEyVcVZVp9uu
MnrR9GEaeplzMcv5VuF/kg/5IAcxDH1ahJmfeEnI6A1SxFauxVGeMCCNds7KJsbc
OHtuMFfJ0ix6jZC9T0eD/IKqkcG/2+pZVoc1m0g8VbK8wHAkXoUqw9JZCwt2rnjA
+3+pLpelMHC6G0U7sMJndlcPxgKauQF9CIJW/9oJFwIgcKmnMdTrTcR3eI10wm+l
CpfXZNzyrwttCDfUfsZ/dHV8iqcR64o2PiEbYGOyGyRFWGd4IjQHZDhgJhsltuzH
6IdvtU3OpKu6f8rsEpEywmxgdLitSkNzMipRy+tqSE9hMRBIGX8asgpVLSu2okX4
zGw8Nz3GSTVBlfIRYsakAXtNqUbIMGNpfZQBGFb8ai6dGW+Z5Ct8dReIM9l/SwcZ
UI6fa5QRouEnqUDbvaH12OnFXTtA+6jsKTubSdTOyzz8lR4Bx2YudaXD+3I4gpRR
DP5pNUW4D5PPBUw5EYgzsuPWq3EDFGE7nnv3QgeQwydyeUHk5IgXMdIZG6V5l8pp
lvR1FYWdbsQoTk7CPtLGqEqZx9VpOUoh2u3cYhvtF+vAksc0NznmBcnB1QJX0czS
oimIesQ2JyrzFwFLWUr4N/nSOTR+IJeEyfx07q0JwmELW3OT0dZsY53pKw8yfwK2
Ee1HrvFfhY17WhoVau7FsZWouSdnjGSbTGlCO4+wC3ehHH5hgT5S2zG8xtsb7hrz
RFpO3XF+s+8xJk2ZdS11GntZ1iwTErgRHWevw3TyWsMKd2chg6iAGx0aHlsfjKpV
v9igABRzA0dh2N+xdIKEHrT94SR/P6r0BXhNagKU4ziNyD7JbMUxTnpx1Wi6a2Kg
spz4IRyWkkkJvrEMKLvDwBuXd0zGVbRCbt3ZScBrY5zs03ULh64wyBqq31fYfp+F
jlYX+VPgRpCuFdaJuaBSA9ZEF6xCeeqL9CYtug4CbVPGb86M335jbhsxhBr4JVGn
EakqvVkiAcV0Zoex3/hG/Y5OaVhknBNa7el4xnYDfndnRaXqMNFhdIwjSCwerjLG
J+UmLwfME2GpsfXhRyR+QYjE0VxYwnJLz4zJUprpk60wMw3wEBXQSpcDC5aijSOf
GC4jTAyblN4LB93zb4hhEx/MnRhAWOSWWMzHdUZrv1TRbt76c+LI0lKwYmcgR1YB
giJEG4gkA4iDDTb/8UlzHGGDodGD4J6uPwfDfnmxzoGUEMFRqx63At2rHUE2mKLA
gpp9tpsudOrL2C/HIbGxyefxQaWVodyU+iqPWeBSck/xZvGWIyG9xOUCyggYmUGL
Dz2z+Ss9dx7CQFr4wNgIiAFFbvpiWehuZS9uFXxqbrxdYNeD1pv9vvEoIx7z5IfN
Mk78vT/JPUP8OZiV+sA4aFSZkTZ0BpSGWi4V8+t/Jmg4yzysscJJxguUowYGGchk
Kp/UCFr1ipdY7qjS77ok7QKuyRUdQM8aEBneIpthUoPYTUVaIulqNANTaUk31Jxq
Y23L1ETficJhSpzlWRG61UAICP4a/AjAiqSI/XJSeGf38e82q+H2eJR1o2R/hN4Q
h6ShR3b9kJA+YIzGLpgad/MqD0SzkPMrCOW6YxiwDjY1qZtKkOtdKcKA4INC/KvT
h7vUhtkKrGhean/9A8IyN+NAcxa9OaEEUcd0FIjHuu+2mr6nvf1t+HafOyEWV0R2
23kaRaLmBvEhxTxy3fGtP3rLXfRrJaowh9tLfzrceilIR2hBORaLgA7MozjJ2Nj1
UCUjMsQYeGbPph+/IYwciCjILCiI6uzJG08d6UeNyAvI1cXbu+D7fnxqb+QyjBgN
rxobdNsYlWBrbEhCJ4pszdxjfWWG4amH+UjO8YsXCbaJHf0kmkeU2imKe73cL1AL
SReuTimmrDo0f+3+zNifulHrntTEFfUes77+6jBzgjSSGO//q79aG8gfOZYIDLju
eMRpQEpOcVyq+9MizJs+T5wzLRHBsRSEIfbZ+n7/VJ9J0vmpH9cGQL4CpmmPvcL6
vpURWq9BBW8aJin9GTxddvpK/GqqMhsoNdmM0CB0ll42iq10BN2WOk6ejb0BLEWo
Oe9RyJHX8nDlk9c/ZKO7nOcXDM1759/KIJvr/HYfofv7EEwJEJjh9cHbuYUH3JJF
f+6VNGuCh4sHU5mKHBAPfSdA3BJI51ptfsOGEof6o99KvXV71Y0xugQqdJrHdoc0
E252satcqrljugm+mhhwlfAJ3fot+nutoa/vuzKspXv3v73joNbcMEDtLKh77yjM
p9Df27YeRuL+wLBB9J4D61NZ2vx3ls19KnShIVg/7ClySCmyf3yyOAEi5Cfv3AIb
x+d/gy9aDCxD3bdEzPRtynBuPKaNalbTJyLlWRtf+tubeh5j5uErVOd3kFSr63Et
YJRN65gC1hokjIy3q0ERIaHTNfzOpluAgo4mJQgFKI7NUbwpdHusjTQ5bZFOjhhP
gqCg0Osi90lp0aFNVmUj8TfPz5TRLQHcLZovYC8JLhu4v2lH24oteUl5ILESLUFS
pdWKFMGG9wZII/9O+hFAK+L/VMQLavC+tNVJWU5ARcqcL+O1BRwDYmrTAMfakPh0
RKUUzwfvjdwQ0svjgI1PbHMu5mtK+cYjNL+r9qemwjNWFRF8rTcm/3JVUlfyBspW
yJRgCcRMia5HrsWFYLzoj/4Q7lI5dqoxPGEOJcmgzQFy9UdWO8kU3uNSwtXZiZS1
iBRZgOKzV30fDfQT/3nzp/D6yvqD/1u1ZEITDdah9vmjDY9WFd1Si4Navd1SIppk
85c6Rnlz9ZRzR91WSQozLKA0n4HQM8m6932kByvjoRkanppKqqJMIz/fO4s1t/eF
LC0/Wa2hhU7qGnMKfbgKYroaxOTgidJrTTMLHlqXGn/3Xx2CaAFoBpWKqUl9bZXm
IKXVzFh+JcnfmDbO+4eMkfmRwT+ZoGhFQkVE8irI9WiDac+GKhgm/HQyLXd2e3/p
mSWkgdavwYx1m9FIu/1iT+TKO9L+Y/v7Mkh3awqbwcyPm18YYRJUlm6JYD+li13J
bTAMYU2cwqiGkXGpx+rh9n1bhwzl4YqF0LAQWkUtjp6R0X7dvJjFEoNroAx46yxy
canfulVfCbmakdktfKPxf5r3OBS3UeZjt6+BMzHbPqXhw3nkro56k+6yrm1CS9ri
Tp5GC4rT3FWVmm3TwAFigCX/Bk04As+Iv+HZiLjXb3pcG53wxGc4aSJGJXPNzeuv
gSG7I1KF0qKJI85iLrFzio9FMp2VeiUg6t98oB0eb26c+XCQQBCWFJqHQSSqOWj5
6uvbToPzloD5CiHK+tmLK/MxXLUU2DRNgeaGRFYe2CquEyTxVMvxMBQSOcZ55Dzp
dfFkbzfyQZ0f1g/i/uu8E4mkd6zOwXsaDg/tvuIAZy3adDtmdawLNmK8LTVmIDpf
GLEL9AWPCFVYfmugIiI9oRlyaaKruA6Bny5/6WvBPNDFSl3wLeuVW4PVkqNfGMBX
BIRX3KBD+AhAr+TvYRZ8rLeLanZo5vP2eokZPRc7f3RqI5U9ZeVO2vvW3Nm8G90c
z99Y7cWyRks3ZB6p/Z5ZPFopq6ov2asUUBjycejDjHg/pMSw09pGRUKrNmPt6FWK
TOkgTYtQq5BuVG8pAx7IFItVrx6x6I5sxMgEr8Hzo/Kqk6IB2tHLaj8WGf56DnmV
hE3B5imARttUT7kTWBPYHK0tDQIhGRWERAqfU3pmG3sk5+dcacnp3zhfe8CHVGIi
dzrPN6PzTEtbzXbBYJXY0aM1ftzSiKG7OKp6GWubLN+3sij9TdvBBTqjCRWBRCo9
Ch8Aqy+qxQFtM9lHGAKQKuADTbt7FYvsdaZCJTVfROhacAXeEdbVHfL0hv6RxZCX
ZB8rw0TDvgTLdlgUcQuIt0fU7vfsMvBsxvGOFIkptB9qyaiWd51bQzi2MTdVz1Pb
xzVb+U3UVJlqKYAZWMvLNgR9coEODepipu7Sx4Kxrdoaj+EahX6BUAXZAUmJceq4
ELscn7NJ6z8U9P+wd0N2y4GWBr/TxJ3ZqXEXjvYy17LV7jgd2pto9VI/J0zfVRUU
wIxVVJh8k8/wyLEwqLxqOz5R4PZVSBw24ILdfbsJXBAcupVrlkGALP7KdV/Ftok0
VXMlXNJBxEgBTESV29eK+6Xg8RgTwWXtH3JWW1G0L52Hi1JjAGIicFSy7THFphDA
MX4bLLB0FcuBZeJOABI1CJn90bYrBL7NilPFqsSoc6VCGORvJaQuBxX0bAW/4Jfx
AsQf2jmZUy59bihrhPy/pMAoKo95ggHnuh1y9n5EZWhpTCXzpNx0z7oPOQGkDoDG
62ldmgJ47+TaOdaRZGF4FYRa7UZfeBPb0GTbxxsOaf4UVirr/pD6OUNLkDlL9TOa
nASk5raPg89yGxG4dyK0A0/fDDOfSHpqKMb+DeTDL+mqYFxYozTKD120gSfWrPzx
/DiBZ3sBV07QZmp3x02EaBjcXg+J0G0S0On6HRhETbh8bGoVGltYwaZqt0aGwG06
lkX33GhN9JBDO6h+Q1II9qgJoIdx/MMXzly90vRdiyLDkngmLLfLOtBM3oNFEAV+
zyAo6drAKcVwdEJvgC7AZSWCwm3a/VWqWv2RzZScpU9iR4h56wbM8TIUlFRrZhee
dtvv50//ZYmRvArGPUkgPmSqQNobmFGC8YPT+Yf+JKIDpt4JghD9/zUIuN+aBuKr
Nxw7S4936cnKUVtEMqmrNB2zUJCUHH6b2G9R/2aTMuZPmVMYg10j0Das8+5IzSXD
PsMj2fNf3i6CzW/ymaZ2EndCutXB67+27JIdR+7v92Q8QQYkhh/sa+3z7HXSrf0a
ljiA7KKa/hR0PIupFErSl4ccm/b+MGTZwiqC5CywIuVNa+bks36DVaWsHrMMkwGM
/lQN5H9dJ0dEo0nVc3TAIp0DtHi0rSK6zctR41sA5lurn9kx9kLx/nRxPs4UCeQa
sqyWjn/0xNIwlgOi5F7hhVWKC7QcDfuYge2ntNvQ0nhQj9mPKw6Z1NekXdbVVlFG
cG2P5NOuVfioM5ymicMkykH9IpVQeqpIqwfM35yDLdGOobr/zWAyN/YkO0j27z/K
k+DoJirkgSnpDI0SVhTjpjtRFEhfkobsDWG0Xww2A/P901LK3IBPgLSUtZU2SppO
ytAqmEHIFdQPhuv+Z0jYrT2glBkKazIcm3nK4i00YjDbF3WBhtack8dyK4CNDpc0
7gt3oq4rVFlKwY3c0mpE2bQ8uqe59cZD5owjAUNXvlJ8E+z1rqzZAVKc589XYz9J
+je80KSGhfJy0wM95+RbsiM5modWhHy5n+amE/AEIIg/IVqlON5VW1atLLnkutHL
uxXRzdCuAq4xv4y+XJxj/bm0VKm8/lsW9jOlUP46fpyGHbrGC/RK4Un7L8O46CRB
peYLMSTCtZNdokzpc0hzR+Ghaqbr/8GnUSSph5aRzAS0bsAal9Xy+7rO6tcVXsqQ
6GNSasdQc98MT4F+7zaSdFVWOT4k3pHnHpXEJGVXUaSKikZiX6FyP+vzEsUVaI7d
Q8+9DctuZ6NT90PIYZdFhw0D+cSUVFhL5e8RSzo8N3drff425xQ7T8pnnFOKqVpN
GCfYrJJYcfPkHLPM0N595MCuhW4hwUNaRjQ+XVywHXDxT+03lBTEC80mK0HP/KMQ
PXaWYbcxeyXEuNT9KCr63cMXWDdn9Z48oQJ3YaBAQ5NRsMMPm4hu1iY6nsDgijfQ
ek0BdYcIMFL/SImHAvI/vMUh3i51IFU99KXk141MQQqTkR73vN82Q9Ew6OmQAP25
dtSy3HC6Gksl5YBQbqXAKPyGWTEwkSB4RdhntZrJc3n3DtmSihi8O/cMnrOUJNXI
j0SdHKC0VIFnSSYf2W1zKH73aiEOvO2KaUohzWsxu9iBmyl0AGDBK9DNRbjfp0II
5SIhYX/J10duN8nUHTusQITjs7ANPba1VXXNQg+Cik0+A8ShzUUIoJuaGZJXCscS
aTyPYQnTwHRRCKlR2tY/E3R3809GirtsrBH5/FsP0l6wDfywN2iw9saOSwwTmZdz
RJ1VCFJ0VB5F/SgBCxVsMhayHQVfAE4El8usjT/TvPBK7MidbXp7iq55/omMancw
16PCTzancw2LdyBFDVKQGwb1kqAxilIhehwGnVIVreZi2BGGRNN6CkguRx+68PMY
nIinCcE3B4e7WqqyCuE6ua3bEhy/4+krheg2QdVfnBWIrIuEWzQxZEgEPjLCvxLY
YASgLis699xqPumFdIzR+f73tyQh9t4vEL/Dh9OZRczUK9Y+lEclerWyylEwxNYM
tUQfmFV8Xm6Uj0YGA+zCRaV2kaGonHEjso/JuV75QBgtjevj4/nvKPSVEL5uG+2f
zswGYLsdTHuOsqqES83DKAV7SV8oTh3JwcgTnn5XfK73p+CvxzzYSqF1U/iRjTqH
4LveNOab3dukeuevUfKfuNINCv3S/H0uy561BWVaMJLvIvLZgNgN0fK2gTYTMJQv
W5PMZM6kG28dGuzb/mr9bsY0ZVcqd8DfyGNo087toY4yshSUKzgYNeDTohkM0Hy/
kZZxWB6Qc6fd3ILVZgGQFZIN1HC0Ti4/WYC3FgtDrCT6VHQGOuu1jkPLLTD6tvkj
IN7rRUemrzMQxK01s6yvERRNjwN8TMwl9MztE023Uf7XK3GAG6/aAWYPSVTwI/jp
7P8C9t8vJEPyWe5vUzDKklyoyoctnkJ8J62Am2mwpyP1UopuBeB9PgJPlhr5zedw
7OoBfFgLEpQZ6N0sSHxCdDvBpXUPEuaxX9PLZcMok5oTIygUB0OUP9eCOlIFItuh
9REFK6cG36AKHnss5gyZdhHpFEqbByJUGTYYkcuSBrVSVTlNxVRQWavBCSNwTTLA
i951gzdhmQNbuZsSPPlp7CjeHo53p2/tu8NfrPEp67FVGvMrtdr6fPyDbNGHY5K1
U6HG7fXLl0kZCtiPGZ9P2aHUZ2yv1vukOvg2FUXhBlCASaqTjj98V3aUu07x+4oe
q4foeXqDe+8h6WM7GvgTervTpsuRj1utcgvtBsGUPyMhz4rFP9oS5Om3Z2+sSRDn
gIxvlndpb+S0FvoIUcIWY3i+Kg3DltNB/5Xw2lloqM6mgsgQvr9FEhhO1j9Acppk
G7+gMa1Qgnc+K06GS60eQ04Ug+rz992GtXFZEC84m8MV5e2iLh0LDNuEJCtqMUb2
jhALML7WltplivRD86adig8mlGwkbzDVTf62yb+dloXlBuQ8r1IH4nU3T4pj9gN2
O9XYKIvsiuCZoR4fYo/QmMhu7eQFGtw+oT7GgK+uCvgxZovWOZCpzQJ2I1T7o/HC
kjzG6gdZQsocT63Rlv2jWctM1ZAqDyGpzi3Dlcf1wOlpEPR8uP4nk2bR81RuAsTK
GgDRyZzsVObAXC8nAMEJNV8bWED7/RERdfOkA1FciFAWxI8uHt9J66Qu/nTEHxFA
n0fVv4JxHrVqrKz8ODA3kafAZqj5UfqoCiZPmqTVMwv6nmt5+APzXHdQxwACXp0D
pd9VlTCca2XwAQNZpPopB3UDZdb8PZSHWdEX9l2vMoTlSdoeZsNSeWu2bIQWoc8s
DIkQdf0vsKqnl19jou9EAUW2zJA2AYbnzLqXrBptJqc2sv5YwwvtGDJHr3NqCqYe
nrfomTnS6MO1Ed4yRbf4XZiwh1UUi97PAsMX09DfRQDf7qh6rUfgCOzsV+rVjnie
pOExuxkYWlph4fBAXDsgIDuOePANXwrGQyBFb6C5L/11txJXi0j0bgEw4LgRfF9A
zIdcyZyojv6JI8X1UIIqqrWLAo5L6PiSk1nDDbngZfM39al1WUAycpUPxINA9fLX
VCoGYlb4ESFW4g/huQb2k9nXF6jCKNsA+OWxKJBEBqr6Ojy4R315MHdKCb+g8bjV
wdvejHc4Iej8NWbwMPP5J+hl22oJ4jUXc1wgIG/Q+HfoPMll1M8DubCewjie7BsM
agXjQQQH3hOz2Yjcl7bQ7xUlCBXHecQpjmyYjEl5AskOSmQFCq5/SUdbJXcIelna
C0tXVgBAEIKbIlMnpQXmi4wJduegzV6mzehMwYqfxy5TIZlVE4od/akijNhi57Db
1/7OzJAOkZuQFFEKtxAfAQrZOoDa09iJdQqnRU4MP2X3sEWqlQRcM4NA4mrURTml
y/4xuY0EyDkiH6k8GZ1l+m8Y+UyY02Oge8hyjfRrytlNgMErzqg4pkGpFKqg6JwJ
T8i34KRz0U5ATuEwKHeXXV+B6ddcu20+2oXoMO387xGY0n464IR8c0m0SM4BhTA4
Owki4xcAtEglWGY5t06YmM3gUQQoKqKUsuzLVSlLvzr+y20HiKFW+FgvifjGRYx0
UrO8FOEnhyd7vD4ZI91KaUGA2GSpPWWTaQKop3JH9U0nDJ01GO6V1v/aJz3nEe/y
4ogfBcyPGU7pFQyRweAyTuBwxD2mCtiKUoBe4E4E2+xY/5vTbxHJudxP621fmdHJ
Opn2ALXCxTfUYM8tDKvzGg//vJt8AcV+pNg8eWcjqmO5Ywff7RLoTVSwXgOK/f/L
u3bRPskqPIxtMhLXZQoaCymAWfwB+vN1NjdX7u/NXv5x4DhdftFnVu29GSGADawQ
8eMl1ijI6Z1xD33l5GO7yCLURDRMnM+kyxn9rT0ey1nwUAyVjzzwFUYZPLx7HC+n
OpRT/8ATHKAG8cBp8yu4rijRbZDV2kr1BPhNvF4b+lhxooipT4ou0pwqvo7IB41N
MVCEa7zuIJIJfPVKuIh8Jf2HTaDk3C36d6PclJ1+7ureUckqhy3zP+fyfdWu9aBM
RomBwZom1KCjJ75LaluBvuJ+4ZjTiHfN4txVoxTEBKNuhbSkGTDZkn3312yBH3ut
653AYRXPo2LP7rjsmKYo/KCvYk48BkVtS7HnGxqXQar/2nLOhnkIBdxxZ5kvVO5J
+SyDY4OSYHCCgnnEp7C9Q/w9sVrFnho4pRZy1ZDAfGbX/Uk98PIWCRExxfnX27JR
IFCWK7A0IBDU6I9tWTyUQ0VK92cs8APflfyb2/UXkJSBT4akhfwYMiH4SQ4YF+dY
WrdIlX44TRLOTQtb6ak4vrbAVPbcwSmWKQ1KFQcZUlcsycAwl3bsM6A+thA9DnJX
krRmOdyGIH6gSrkvPxHkmugoYQ83F+aOPidihsdBFAgWnZHn9KmmzOLHAff43OtD
XjLoBTx1LjiVT4MQHx9qDREL4pk0Dr2lgNK334i0NylsWNeS+ikkNCq+UzaL4iRo
w1fxTof5h2muPLqxd611r+dV7saAveb7UT9U20T5iytai2zt27zTHuTgJmf7UaOY
NcNeSHe6ooFqxy9UVrWgip6jP5eYQQEF383yqI+DAxCqJvhyAej8lpqZZdAmKWb4
a+v4cIOjQXW9YKUFbohyN8BeWTGtc8iaFE31n6fV1aAnq2YDngXGbdUBFUZygYg5
y63mTCINQXQzq7StPq582EGE3R4aP0cxf5KJeC+BBYImbGgQzhq9SIWdOcywjFv6
TwrPeqb57Z5EwW2hVc1rOr9WNJzVx8eTUHJfRZ7/SYN7I+8cu6D2rjcThvyuuBdt
hsMYDIXFYL3ZO+zpw//VQ42ujpbHxvG7S+/+cGuWB3TZ+1hXpY8zyIIIZHTE2jVE
dhF21frWUOComVjXtUMW5QAW/dVDJjf4JzNZ3nzmEcCCD5CY+Plh386ULRjvI99s
BaOJ3Ah3gSH6m1uq3wKJW/5J9IQY8NPs3a+9UtD9Z8lSKlc0NR53g/3R8pRe9ALZ
REY3sTX5meKZ0OuBQr8IFv9xz6PxUyIzxyZWJoa5SbJmy8n9hsnRyWC3zUgcG0q/
wj0PN354qMQeQrGTJ+a2tr+CfgdkszK7R9JEuKp6R4Wsl/uHMXY8c2eS5c4RDDIe
0U9aqFPv3zw0sVq7vjqENdIKJQ8/HXFkKqQYUuMcESKM0nEcWtWorvqWUnwrG3hF
R4SlpzuQZqFEnbWr1ad6k5zEyQMMLxLRgxmvbunTiv4QQ+q2GOa41huB9BOkr/Qk
GanP7ek1bEnHeXlGZb0jRRgDlt6h8nEeu6THof0PV4z0xFtBdTRoKkPCeKa3e1CT
KwkvxljrPTJAkZfNHay6YPFvYmww22guEs8hgcoN/kO9fJ3DfQkGJwcxlPHXdV7G
ONC4dCEWPydLpkUcAzItSxTj5OmcVp2a6poRvQCJmE0xokWcRKjrg63r1nd1lwFv
cJ2515uhsNBFXFLiWgyXWzBmniur0YEuNzy4szUJhKRZW7ng7Xd/o7/0+/TOgFUK
9BIe/jumWyIiJ7qY0m+GG4lk+5hDPWgWC64cy6/BzcoPTzWT5myc6JpVmFkLCrgq
0aQuGSqgspUE0zNnnopJ+D75FlMxDLCPchugcAehIjSUUPURVC9fViMfuI630Vd5
WN+/BnbcwaJj6ywnkO9Ms38nhiXhulejN23uUfaqPeOHoWpMX5L6hMHSR39N+EvJ
TS8lPMPChwgOpU8Tm0F7rAbszBdFxuEzkNo2E6xENyBNDWOvkjOpfZ6hLNuUKkrE
FML0ArwZCASNvAqG98T3sT+6VODc48mfqZtr3j2vDky7rB1E4FY4G4ZliasNZKvs
AABiAwPGr0kbdlRbLRZtFeCTbbRhU/T1or7TBQWOVhN0oLn8NReRMUluytzxhEyq
ib3q+/bsCZCuoTd21z0NU1lBPg4t/MBpIAkJtR/8gihL/pT1vS1Ie/flR+hsUukl
PA0tOnm+E3cTry/Z7Y/WHdjjRdrXPF/CdSLyV3CFyuU0C+Q4Do3iaQrshRow2Orx
4hnYyTW/HKtrHrbT7CzbzJi3PwzGgov+nCLruxPfNb6eucKK4Veen2ik7uoIcn7j
J9SWwPpNBDUN3tSN3HK0SS57p/1WGpyf87u89SwOVvAwxUWogGXY/zYoJfeTJgHC
+M7B9U1R0/xRUq+Nafs9n3Hs80wcQhDnjv3IGrPQYGwQc/+OaUwlXKHJQbzv6lUT
ilyVpa76ikwOb52vkYkgCTwZ0blLUR4kGEnH0UDxMjVvS94Y2WjrKlcVmzfoh8Xh
6hlKk3TIynjx5Z+LzuVWCzk36JAR+ytrsf3FeOZRPAK6VrFNSalHYSJlv0MBo1V/
wFkiNkgGASkFLQEPQ9tjUtCIUHy9f9x1y1RBVAPyI67XcmwswxxXo9Jd60YhPPZr
KA1TeHUeAvgECRP9piGXKQqrMXVGcrVtY3wPLk7y233vz0Qa4dZHKmUcMkWs9jK4
veAkCwdp6LdOjra7xaYSSSTS6p+Ig0APbAu4PloJL5zBaXxOGjYGxCKZP61p3YBZ
Du0KXZqHOHvdF09hHfCj/VTbzQ7B9yhcN/ejuzF5hkbt0wXY2wgbunY+EP4dLYNj
BC2M39jFZROzxy/Suz2OrOjg2E5Zde5M4JMVGd9UJRXzF2KK6UI70Tr++ctj7eDd
k9Z9LoJ4+khem/PzCObOjVTjgCD27BgCP/7eVtnChnBG0wUN6QQ67zo39UPW6QP8
HBVz14p4CCPxhrfk5cA5DtXj3hk0a/Y6XW3M237WtmgoyI2LyeKnEw9UOWtgO/cD
bwn/fQNkPbYybyPqiD3nOTfEBwqG8J2LOa10uvc/vHshRoVKI8/nEwr9Y3ygyKYO
4lvJJr0dP3/T1GUYI2wVHO174Cqq1illdUZfMLPgSAASwb83c4ghFAE6pMWeBPMK
3cAdM5es4yzOgUt5/b2VIquNfhyZF9skhzTFM9plYuxUWkr9bs05pviJMSt6BjpM
USrkpksx/bpjwr8g9xIyb2exVL5TaEDK+i4KeRJsRc/IwmiNAT2nu8XGXggcMBUx
ratfD/DK0XM+Ns2W+eveq16VoAve4f2Xf4w5akKwUKwT9y4kxJID8dIdYjpH82qI
SdyTHnyqqtElz6t3jDs/H2QsthsSodGAqKs9ApDv0eyAS3LJaBylEydiGjFqbyQU
82MkEcZhVCUbD9zxwwlZGVNTvNKxxgijLxZwnWmC+9yINUkz3iQd4E/hAVapB8oH
uJ48CYOB4YoYC4Rjy7t4C4H/WeMbmTFkJIsYT63bYe0u4H8DhXGOIyCkwbMAnys+
RoJFf3G819q6YM0spnYC4uy6L3Ro/SOKxnPRS4kaeubTohMJx5Q3vIJwhReEM7sJ
DQ4tCC+NeqNOR3r9z7+YWULrJ/+xgCU/XJmz+bgrWfsQxUKYZVONS2Tw8J6p8DHY
6/F286qjfYAoX9QaYrFeCZ0utRRPXVAb/+21hZ5JkUGdXXfQs7SBod+ecUrtupig
oBH0y5fjm0TiJG1kp3YylJSvBqtUtp/2nIBMn9eI2u5blkG+chQTTEU5E8JRa42c
LWKbMvljHl5U3dyP6Yr8iS7bTRkEIs4OPiN9KxeWJbR+NKs3/n49ByCN8V/qgqRI
Z3hohZwhyHeXPvhfeGw9p7CjWklVbbnba6rxkuh8Ccq3WhOgGjKatYizYPujsKBX
8yCvp83FUsjcsM4l/8YBycxKETBqXUlymzGw5LV1ipcqRiGT0Vzfy9Sr2UNr6O08
FEAKIESy16ZcSHE7Bvx7wzZ7Pd4mwBDR6XjaEueW3KMMBYiVz4xBrOCAKaJp8maz
4A/VmkcN6aSKef3/FqKYv1PBgyE7yoh345Tdak90ITGtqcfAM+vM393e+KPBBKVZ
e5zgaoq4G1D7qYnq7cNG9UIZIqIi+/EeYwj7cW9it2p+hTgUSltmmCpTDVWBnyGS
D/KgP/Hu5AT3rV4Yt3S02AngAsp1MeucK8QSlZkOcv3d/niF04b9JHy5ox5jU8ec
4KhuKfvlKGPMlduaW6QYUoR0p6HJYyG+3rYFX7wN3tGv+NLrkvtnYc5X3Hr2VgVe
hMDIr9QM5DgaJAnQglhOckDFp/ZzOuCWQG7nN2HMGbzb00KH7Gxr78FzcPSiEBY0
S+A3FSiTbTDV7q2bEn/cekcx/OOwE0aI4Qu2a/2JLPvsSZn/XJxvY/c93/EaK45b
jlyQ62jjd4vRIybOhRlY50BBKWU9UFJedN1vyKGBpHAePPSS6tywZeBNWlwfcLAq
K+wrdjt1d/lZtEjL19WyDXvJOciYLyyekeLYFC5GHUDRUxSboJZx3SIlp+1VQz7A
VBPC1N76+1jMLHlW2fUf72NBdHClLOEOeJOVHBKvPVmsmMXPcvjU+kPtICL/alMj
qN/uqdgKL8HwRYDDnbgOwgnp23ebaaK4PpaVKSHKRUx3A5cODaicCBZJBd58p/tZ
UB320qFRiHoUqwYBjZOd5t1lrCo0Mi4XzH5X4vbMdNgswUOQR17qCbAb8OsAawxp
5GMfMzuYYzoMp042FgI0PzRDFxVKfwvyugo4nEllk5LSRNe9uEMO9FCO0VREktni
g70WWz4eDTViF2//MOvYfVVWsi3RYQwP91QV0cO2B5t6veM28F+HkFc2l9btR0oZ
QRuviAkDs3Q2F2sFvsJyWHrZh9o92ngT/Goh2rxL9T3lKGzLyMrMn46BN43qj9JQ
a1k0N+eh492UKsWGCtM4JzNsASpi0Vyl1pG8LvZisghdU5w5DN9MWX25Ho35NtO1
LfYbcRoH/H88ap2iJJfzID2jqt1eZt4viTrzDM+wMnDp/K0NZGgi+q2lEIpUOYdF
A1X17hsuvr0js4el3hmpiV1FDHFvB2jlLYMkNQGKg/atOVVgoTDlxpLb6E88P1Z9
OCU4/ha/+dtIqATPUvl0JdOCjXsW03zfCCtIHxHP8YD2ZvTtW7SxxFnmy37+MZb5
BMBSMOXvTNPthgYUy2inFSQFPPQ5Q7R65V/4H73hHUjG5e3QP3v67oUAJ678zNQu
FyiR6FmjXFR0Z2DQhXBRfFC/GMFkeEDuInNvo2pv90/pzzbjNwkAGhQ7TJ2BUFpv
KljBk9jtFp6+5iniHQg6RLCFI0zEkB3hiUyIaFUYL9JoZGY7yIwcu2Dh4HWPZMX4
AUUgsbRoAQCDVkxvWFLTyRg0kNkiy566oj6XLlHHAxg+yJ0chCiuzuSpHbdTEcpx
PDGL/TrgmuGpDlAnbZyZx5erO2QtcaoD3bGKkuctbk0UACMgpqCYIPcjjbhv0Cxb
QgAjC12XIRajjeucYPpwYVOlls54G/YEmRtj1zrfLe6kWmWJUsifK/cX7sUuHvd7
IYU1jNlTcesKefFIseCchbAxOBlA/E+xt7gjBqFMPotr6VRbm2bAeyc7FhDosUw6
EZZHQaBZy3szcW2PS6+xjgBpOfDw1oniqz+e25+sQv1s8myDIf1DkrFjBAu7E78G
pxDucNw01jNGjmBHtyBk5ax32CgjlGSjLmKb2CLIGAEXLLWACeXKYDQY/I9wwpbl
5AvHoqltjVKLAqN7/3r6s4bbD9bdbjGM7Ozy93HfZyGWOVx2/5M2NVX0tO5B0Jd5
sR0uQyyNn5czhaOFIFVmaovxu3xoH4JDqEfLp47SGxq/KXw8buquITaJqpzESbUZ
8c//4vKCM7Hvc7xoRFEKHS97dJNkqimDotiMjyoc1T1jN/79BwVnMi0e8iVTPnhK
0xEzsxqn4TaRvapaqDhi+bSsW47+jJ/yDC4YfJQtdppioJnzBIeZgrHSzd+AtLLN
R/hAB8rlQx7AWtR+HMGyRA6vIWeGIZoitUql7PmJxAfLtbnJ9tW4Nw1hIYWy4wst
WG84WH2gQW+FX51qEUohbqVbGkkYB2MaJV0u1nQJQ30e/a7GO2LJIU+zYfYBtu5u
SV8Vcx9ouWqd/jVqexgezl0NJmbiQZos/iyeXvzO/PG423Or/vuUxGFOdDwjLML9
kiIPItmGxmGimyWAkjrQO8XPNfawfg1ObAd6F/e/fU1PaWrVK00+zg8tzbq98k+L
cu09juFcbaGpXeXhurHxJdPbeWcoqoCxCmiK4qzhylRWzZzDmww0unfcyZjsdkbi
wHWqzXmM8IgaLYQbinZ7kmtsS+HVyDfRNihXao5UiIyr+ZPeJhvI7zAimwo0S8/l
Q0Oshw0ACZesAIYDJbkKaWsYPWNG/IHZlHNZ3SUhXINRSGZ/VSK+LX4OS0KM37vU
N1DxwDrRXY7q/yxFPCcwEwtr6bNSMsYTkXXyPtwiTK0A2V5pMJWPtEMwAQqUb/OZ
dm5xWr/6SL9UwmdGdwA7eSMMxrga8h+Es03OZCqEVKiOm/FOmcOMijDle8fQoK2Y
waF2mWKQ5TG8PF0RPdwohIJYVNHtKpbGDt8bf25YyMHgoLCdcLWbg1AMCmCsSOwi
bWSPzgfbro1GZLBxR28Ykh1eDdydY+S2e24HsEiwhZngJmliMXOjPHYVtsIfwMNL
wTsCwOo3zblKj5W10Js8ZNvni7HCmh5ilcPeO1OgwC2gnQI2SnPydxRtOt9GFiOl
UQFs6rWwRbyH/63zXa5PPs87Ju+tejyVcKCtNRFayCotwcRNblBAK8rY7jsV5A6N
St1EsNseoC9VOQuI58nZuA4bXB/5rZf1rkc+g7jAETKn3fS+sQ4+5vhjQXTRZqcR
/OGDv2t0ZM4NsrncY7DOfxtPhm2I9AyK4e3xUPziaRuKz1ZWauiR5z0xPYHgxzYy
GqucOK/isIkbMQi4d+DL1B3QjbHHwvMi56BCAalac4CwLgj6EfRLPPXXT68mGdtZ
xkTYp1mJSiFVcm1bUtyTFqhHyWOskbYr1qciApOH7sh1ONdKl6bit+6arcdcr2on
8VnJszrGE0hyh/q0HgiygxHLbskMg95fIyD4AMDIIewrx6aNI8vmhKPuJZ+0kS/f
ieP8ZKjUCG5emApPPjzwvvwyz/nHTYy4IfYa/REwrcWBnAE3MoOs42WMI9a5KX9y
1hzBheklkciAQrgWL4LdppoXoW2m/lsEi1uo0gFo/yjBaL/7/eO05D1k8LfmF73k
M/WaQUgiogVFD7fEpCXi8ETHMXLYojytSR4ixbi3e4rgDN/MhZW5xWx9lGf1B5YG
SydgPQg7AdwnO9gE7UIRrH3QcEjaIdjk40jh1ElQ4jmU9jPzvYk+I5Eumh5q727r
Ikce0fteYs/KfaOvUVc3a5zhuyQ8GJV2kxhbNggCJ3DJzvo30Z86/iP33bPezosQ
he8NKxNd7bbRwvTz9FokJB5D98iuaFVOYfJ8MW0cDep5VmOSGUeTbazrB+VOBe7f
YywbYV44FPqLkg+dZR3JFb+z4I/z/jl746JZHBnOvqVrHVzwp2v87c4G581SJdr9
k38Q2WCkGA0/FS28KDW+BO27qx4dluj5hL/F95ZcDQ9ji1Y++gra2xRtlHo5sG7j
BYkeMFZoyrw/fkGK6bmiKxdebIxNS7w//DILUaoEjKLpQ7UIGbf/72cfdPNKLahL
1z/qezODEJhcCIrTSJk9GcavVB02Qir7nn1JIT5/G5eCs+6FEApK065srDi7n6MN
E0TIjsnAHkwA7AweKS7wCkf3buUu8ow0uFOLUXj8NzpWGA6Zp3WHWGAgUjP3Atco
uUQEWJV6RqogzhgAx/Kj+IduUYZ518DbbPQaxS5F8/8YyKGM7UX3WoPNT62lmJDb
fOL2iEHD2VSHxIJm5k8SgYxz8I4+O1a42kHeHK4mQJ+zlOt/fLrFtauF+RuiDIlQ
lAobmjaM9RUO+Dbi88Wa5RraI8QYEUZinZjEaJUpXdkzldD/i+dxlsHd8/JfTUPo
0aEmdNPpF/nWyW1hQgQuhpRZ0WKfLi7596Q2gU+WrDbVt6akQPptHTI0m4hYa4/Y
nq8v+pW1U7eYOHxLhL4Sx6PbCpJ5IDQ7oU3SqhZy30d3JScaY7lhfwhcUdoqdlPk
MLDFGebbTB3derodcni+O603qcIWmaOMM8/86ZS7BlnjEnSj8wM3OStYlDUQdolM
FXv96oRr8CvIA4UwqqUsBsJ/yOyH0FS4MAcLN6oZCLMa87A8INJwJlG413uKDsjm
phmoFX4EHjBuM6XQ0GsoJRetVTwXCKsOLGr7UUqBn9dP23H2NaRLfR+Hy0zrAisF
rEGl28OrOHvQoij2jaAYDUZICJBxI6uo7AL2Sy+MbP0faW5uZiC/uh7Vx7pIjVYG
WoYDCO+EjwRnu7KRIvQIHPHfGxbrzoYl2kVUXgzHtEfMCsqznDcRYLZS7swbnP7E
jaHFdWVvxjTL9DPoSeRj/YQl4Ld0RmryjdDPndWUqFEcXsduFUrPIpQlmfg9M0X4
wKSPg+D7fE76KyEbLYdFMJDe+Ko85OLwDlB+ab1stgRVQ6Kct4x4ATCmTt5W1bmj
QUdd/DlrUO5K2rNarL1wwfpRKibH7olaHXDXdX2uKjx7z1vjOuTklwq8A8SHD1Gp
wO59tRiV/rm/93XNob9wQHjAZQn0rSeqg5HlO/E7Gxr697wB0jPrWlEb8K0yQ1i1
labrYyMDNiMOKcS45VR3MdG+pnh2jEGE/aCcZwmPa+phIIUS2ysK48XN9uq47FHE
Qyubj/AnnDEP6FpJfAovDUuwTEL9nAolDajpaiSJUKIj7IT++kNBPd9cenxpJho1
d6AQwD3Is+5o8gF2L4smG5GYWhyhg7O3wY6dnOVZKbTlbQ4tnNuOAaYBxesfgnBs
hyBQRGhDZZuccwlFO+T3D1B3VmipZQxQIpW+oYYJneGyPVJNb+L3C55+XmWLT9KK
8n0TKN6uKNajgTpGQGcyy0J8kIIFo3tIhT2timzFTUvRi9GjzIOv5mOypKtN7XFB
EkbxKhJ1VsvmznpyMqz/TQ0gs3C5sRjfw3RWibqVir7JQAUEUXK96bLjZGQUd44H
i1uCiecV5BP1YV9Ag/F8wRVyZfuNbuv81tex5A1367wOd8m3+SmN730/wN0sIX/c
+Dp+LMSxoZ8MWWLWOKlbNwyNppJkVnd3yAD3Ek9sn0MC9d7tfwEuuRkkLjIItVrp
gcf5Bsdr/YKMc1pR9W1G7Gz8FipY/LDHIgxkJEyIHF9Z/F8fGm21N+gNlTsqQjX1
bgarY/lJY7HNvbtf8GlePoEGoPak3AlH+KQDvtq+sr/3L1NiHcGhQAN8TQFAqqMv
EQNK44+ugEOzH9pUv12I5pqVoJsLbnpBynGtusOD/h5fl3xlqb8Y4Ordsg/DkJHk
57lfD6HrE8A1Wu+lP7/v2vvoFmvvuWDTIdNq1lUozzsroLwGlubPfYSHN/ZWMzQ0
/QDkX3vDxAVWc4uYmSWuMOP3ry5YLiqp5ahs/KWDiHNPB0vxTFq+8wZXqI4PUKaw
OQTZ3pDZmDF/83kyZcQY+BsJ6M508+YnB5iinTjES4hHwSiGTOVFviGkC8qkDVRj
gO7PoXXuMRtDQsH6hWWLuykQivXevYKizG2j2Nr4+/fB7TQr0RUYI0SvWaStiY8Q
hILZikDZafsBXZjsQZ9nM4/uEnh3kpCi3O+3Hb2AaBKQiIx0fP7IBp912kUjLwVw
zabk5kfOE4IXDLPagdZ3BnxHNeN43wGM6f1P1K0PvTiTWe5D5Lk0Z6lsdlfkQedm
RPq8j9lwtyPjCaQDNUgu9Eo0FHiTaea0qYlVqXGbs/XMQQJeghkTj+A9HylCv8Lc
HgX4XjyaUlhS1UZKxKC9ietHZzCwjycUMxCkgBCIBn6A1KH0q+sx7s7O6fcL4Au1
EjU9XiEy4qywCxRkOebKn0fzdd5ji/Twh7S9TXgChjJs+Ui44ykqy0swiJKbYlkF
oc4UYTjpt3LZk/N7cznpHL8uh44O1JRWhgaaPFsir6x2JH3TPr6OA5VILziU93oL
GGoxcRkQ4TPZtkh7KH4fWWKwWr63zgLdUky65CZ9idCuX2vp7jKAslkUOTO9Mm0O
uvmDI6QWBewdJ9tyB8m4DQBw/yQXLDD+ovJatvaFXCSXe5ntP0kbiXFOUUmEQc73
4pmfyYoXjfM+oBGKu+4QydPM1tlWMYN7UKa7aXKwn6VpSo/1PqgKD4VeTLEhvMuY
6ne8lR/95hn8TLiP376CPmNBcUPuMeKkcosUM7yRH0pQ4HlblGNLG3i34HBSI1Vc
8xkaGAu3YcbEl8iM1k/xykZwDibE/wGNMuUFkoje0jH+l+zU+kzn63eTB8h8gy1a
V3UtjLKzMDan0uqqIbDL1evu1XQd/ZYs+k77nhafv54O1jfqMGCx8/1GDnxk0yhW
FpLymXsQRufTo3LDywaHyO9li622kD2r7O3qeIZQzVBt9/uJydMFBUICld4UeBQU
1E/xCvznJVRWwptr0roD+8oHcpsGvaHjEkJ0QQ38KK+iOkDZkmIfA8kU6peAJQox
n156mtdsB2nN4OTU8BIoE5g5zdn2d5dmy82iP8oi9NvjLB89mDTkJg0euTn1x39O
E8NYgdoxkVtTFMAdzVIuTZN/ajiczxTS2+JjmjejKd1YQtxSVRUcONh6BAzffBYh
xznECKYWq+ndJ3wzZzX6WS87jXJpSJnOEq/ruwJhLO/jx0k/8e9UgLXOyA1H4QfF
/38c9J81slHifLNbtfK6AKJnYKEANQ24vUeQhTZkZeKl52fLa1VK/tmdGcDRKTNH
SrBWHa7nZN9dQ9g20jNA/YZbmnBhTTJFNPgZU8EBWv8dQFgtyuXv/Wc/rDRjMpLa
ycW6H1/1M4ZaAdRsaxKHXlhCpFZYx/HbnQEvVOZZaIh6fLu9+LoSQrYzqtxxA+1Q
xjABRWNPdVV7CRQnZl1wHQ8/0+B7rcU2qvPQUcwgelVZm85R7JU++0w8RMZTIa3X
Q3250h2v3y/Mmu6MEM7lDb2GNPTnDAkBtt/iXapXDGB0YU3RKMovZJk4/kJ2sz8P
YRJjHsYQIyQzXHzEm42Oqhyw8uQwICf/QdLaYIZddPq7fqEDBYD3ml0p1iAxQ5es
mzaKmwEqOcnSiRtUPpr0yOsVXn+1vLJZbCBdncoPRyle60yXpc9ijp+CBlATKaeO
APezcI2eZij9RjuE9GsuUQ3+Lvr2NEWrw7yjb6CkBNuBQAcrLRtNpr28ZyUutkDy
Fkbqoq73uTshm8CZXHkbUEaMCI/3Rfba9fpuJIN40kvIWxICGfzvipU/6/k9tlqH
2jF8ThsSMkplUZrPRggML43fuUlcPq53wz0nxQiXm0Yg0BwZwir087FK2DbEOSF9
UJHFQv/wteKL2/CIYdDU04eaz5Y4MkYufbSmuSzsatK4gtrMMSEgFG0i+jNe64YT
LMh3TSn/RMc7D5rt9ANMneMteJNyjKY1RNAdnBe6jB/HpJSDcwCjhZMCbFpA74XH
Bkro5zOQ0riuPxyUYF8Idg3OMNa6KTF2pJcdQE+Hd5TtkhPo2VFjfwuhTNtlUuzo
0vMmgM1yr8zyDxNG3Wp0+inC/QbERR8WYel/ZSNk9/U5jTZhtMJiz+gZxflW9A+l
s+QrY+R6s6bWnYwB6eooJES0dsWoFk6G+YCrD2l8klUsCVhqlV3aRhlj7LtzR2jD
PPwaZEQ6DCpqIY1VsxrSV1E/5Fnr1J4Fg9Ws9a9sBok+vnLg9Vvlbr+hOEtDjRrW
KD4kUeCq6BaAm7qND1dODQazPRFMRhYRaipDEvZxfp1cQZRONr+jVos8PzpicDfN
rTz7p8vmpTW0rlK9PhLQJ2SvxeX5PA8g8ivHaF2Icq0rPh+TmrIQsze8d1jh6Ru8
qBvQ9P/fFA+HRzhNKHcjudzG/U/RFg4RfSu9we2EDJP+dehuqQIKK1J2yxwkTKmA
CZz2ea8oMfhKnxkjxLOdv3SNV0pMCyD0dKHTgpUI2uj+QSxH7+D9rkQRsTeWHofD
97Egi0bbpFexknE+FA2kbOhxR0vZfsW1VFZJDRdMMmKbw8zZwF9VqXS03iosy0ZU
6NDpgdZ+C1OSHavaMEAPNM4Zg6090e7xTdNeGAur/AUDhb65evicRC1B2k1uPwv5
aC/a61REU7umPDlu2vfc7dBiV6NrPsvpBuqZT5ZmR4mQUQOMhA/gakvhz7DuZaHT
LRnNNvB5yB8om0gW+9Hhry/XQAcDcxv6MKFiQiY4R3ZNHBaVCQnrlg9m6gI+ZBDp
yiPR89o0iPvse0cxdZMQwLVnj0dbXpB1TTfboR8vhghe99Kj4EMO7seYeaUvAbdb
7p3VSsweEee5rAbKgUkD6NbwiQsMvUzjTtVmg2vAtB8MnH00mCR7uqF0P2DLOb/i
/xhYut34+l2bw4Z6e1rpmICLJJpruBD1rp8Si/kR6wFDZjLH4LgdQuedUi76is/L
Loq38A1nYOwPvM5ycDMpxtMmJ7Y6Xd3GyQ6DaJNOs1lYXVO6nOUWjrLrJXFxjqV8
Bcva38PYr+ykCMlXTj1p/6TWRfInjofACy/prhpwpC7+x7KatIi+HqCL7iITbSim
EjbgEvZGapSM0fl1qRyUHWDzxgutSTs7NH7wLiufPyxyLM27N3ZxE4IObhb11JdU
AWnkopmnVdrhT1yvsTtDaDicJ/BlGARfUCqROH/ilBwbio3jq7pbYoHveprnYvfH
Rmv+hJtury+YcwJ5eL2XDtEMlST1jl+cDYgqzCpqakdgW3v75tFHyfjDJON00zEw
aTCs1LWIhaHr5EiOz8nnZnUPKwibjtdrN7Dy1ZEiuRU1oW7tQ9xhWwx35UwMVJor
h0IlvuOO5N0T8UBnLU9iKjV43FbPgf/m94j85JWwjz6rOJbyhI32Frnhh/8v+c/f
CBAhvdF8eRIiic8GQgSXl4s+CJZmfC4u3MMa7m7ZfhXgIL/gWn/E+2XWUxspBpFh
G9PLeMCT2w65XrvIo3yXDaxt3MyAyOhUgPCPXZVhfn2rLkDNAzAZTYQN68PhzOQg
ivdktmkMnxev0BH8cm+CgnPYxH0Kgl4EkyZHZnN9/ZyySoyQMXlzJrjQQOEg1f7g
PMjXGizgb40uvj1af7Mf1FLsIDSige9oesMN2LwzRcO/IfZ7PnXRPSIxOOgjGsCb
Jmt+eXVniWvWF199pkCz02vJwqdQp/Wpvg2KVYSqDe0SF+kEQstGy/tyV2zwvC12
WsIIJqofWSw9bxwFmGcrnmi++5L1vz6rSIx7lE71+j0YjsgwzdZLlFddKSGVEFvf
2xV4/OOflpHQABPSYuh23VnbeUOHrOLFvq0Yv5fUTbhZeEq+G+P3qn1NWxvqXbc8
U7m5NSsX8SS8IFN6zf1KDTvccsnluwbUqM/fOjpnV0Jl46nmgkRZwnJN71xN8okq
nPjoY635vndHeLKbgB9pAdwvJK03IBvTjgprT16/yYx/+CbWMEFGQcwHj5MgqrXq
lPe9iq28RGNlNOLKXvdObzP79fREZ3LbEPX/ziy/J4j6wA2Th6zZi8XX5owWamKX
8wuy8CQCxbFYwo4uApNQ8dTRD9Pg920ef2+GdMM6WbvKe7UbhYdQWiuUjuBWz4pn
M2gwcN/vuRf9w/S/3hbVoCrk6Q9jx9ZfSwlAFqo8Wd+ovJr3iKZVnOn4J76mk3iJ
bPxtRAFgkw+Wk6PG3ANArL6ojxp0JWnzPZQnCjr2QWN5RRQ8BvUHd9wYuir20NgZ
pIjAp3M7ji2z4iBAx2Clv1tX4IuV2h0uMlvxzOTb4U0wfey0iotBIip2STXWXUWE
4yVcU638H3BR4DM2RyDkfnDktofWIGGMz6gohRVmuhrhoGhyvQk4JEp9jnwKNPTg
K2qAXjVVBAjX/GaTimulQ/+jl8NbIyYl62rhkXYMjJwrKWcH7x8k+mtrkPJdjjpE
J07PPpV67GLhSNNVUhxIAd9/Ww0fdgOnlFPs5gy9X5T9YsW4KSd5RNVxLXNZ+iNm
00EbM6p0TmDdoP6N28M85FlpGR7vUbrzUi9ghtkXMj2YsMgUYhLFu8Op5CkjaHC9
nPFvFPlamS5NPVjSaZ7rVu2G2pwzlMh4FJBEy1Ec4nG3coWJzSVxc54Lk3sSRm27
NBC7CIgLiHxRDy4lbshF1tKo0hiOk3cxbdDpRYnZSVgdqMb/CrA8K1Ez6oXf7KN3
XykkkJjqvx4y/Kav6Jiy1yDPpd/DKVoO+xm5wsx7srWqsrZ2qfa+ejKifZQ+AedM
zFAxN7tJbhCp1f2q9cVNRQM1pnxa9A0q7nfxWE+nJAfTDmRg61DaetvtS6+OOz1d
lczv3Iwsg2EJY9Gk067pj1J7zjTD952EXSYjutVLJyRuEJUgpLXZsg9D5UsL1OZg
iLH77nkyC54K/ww7qjJa7WTafjxKFpwnFtAWngeZBsOEZdn84iPVjj+NPpZZb/Tt
2X37RvTKosnw5roP6HqV2I2ZGdXXeAM0A8U8YmOSefhejh58alNh5xwg1hVSCgnR
/zzaWc5rhFE8HZ/JlrZI4jU1xTykwJT3TN7jPcsn5zGpX+4bOJULKED6OWTzbP8g
/msmZH7HmoH6TluR9frNhF6kJFJWt8HQOk8WQUdeIWhBoyyjB+EIWuuhZgW31TGv
IcsTjLyLhYeAv4MdcEZ2Zq4hhCwXl1+MnurbcI5bIcnM9HKxqrK4eRIFfP6/pv6+
UWh57aX1E5ZckYiqAq0+kjPckwBFLyTY9hi56lDy56JrOjmzQVqJXk0jh5u1bePx
T7O5MncLfQ01/GZ3qoPmUCFMvRh0NrO+3WBhFPkNY2KIEaEgMRf0YtWMANO9EMMS
PVkb5T5XIrlAdle7EH1F/Bzd6F7Z+GQY/1KfxhPgmcrpXH8t33w3Kb7i7bDFGzJm
2FcQ7ECKptN2knLwE3YQW2CeMRkfBLXL/jUeMUI2lHFDY5l6HAIbF5FvhiY/jFgm
zE+tWtof2bxPYUz3XTNy4D0caqR527fR79F8PToKVLzNIb6IkTnmwdFsBIzM1HHm
2JUkgUVtuHoEnunPodlEMb76qF8AQFfM7AUyHfXUB1oTMdWJo43Yg92bqEdNR5w1
ju5VpJG9gD/XCAsM9YY4BvG0MzS2R6k68wyGlE8vt/AK1TZJfL+f3i9GmaFpnqw5
csamzqqeBl3USGXMOKIdj8kcLVJdj/JeuhmwxNZgUd/OSdC3tusozNnmll9MlXuu
Szd0nENI8Bma1p8q2pZ3Qu//hFgBqHypRAVwm+VTUtJgL9XWSFbJ1x0rQw4SWP1i
TaIF6u7xuCALwqugcvqzuugsSeZk8Op9M3D4g09SrfyrK8RDu2a+T7LRGT+/Larf
bdRAkicGTLEUa3cJ5SutRDGo3hmyOsnD4j64jscIq8NSYQzKJR2m2N7MQEE6FXod
Pa8nTAAo12QCk2NzWNDsE4Jj3kvMhLGvnmDoi7Hl0A25Vg/jXw7OzLz5O+I5P4H4
1JOpMMIa4tNKR0NHe0yhquz07A+vt3xeGg+muUSXGYE8n+5EUVp5K0f0T8gpCCWp
f4yikoHdWkwcJSxpuADC0PiqV65YPiGjTynxC1u/Wl62MMkrdpVLatFb+RwdXgJb
vGgV6nbS7Sw4m4S1/iNb0OTjn+HCN06chZPb/LgPsFBKs1z0vNZ/hIBd4rG6jqrq
GM2TSAYMABVUqkED3uhaahom0XnR38IDIZXcj9K8qMLF02gNoRtHMedv76hEr0oD
jh4QbCnipQoH83iFRWcc3bxFCB2K8FmI5qE0/o+3AHG5qFa0hdxJh9Xr7puYiXVT
YncnYkFFgs3PyRcuZDIRjqICLEfO07jUpFiD21T8jCrHrzH02q8KaBz6xhWd1pwq
AqkM2eMVVHQ78hZh6RrqyME7/Bs7pSKaCmw9qlnCCgmy9vFvWvPPpz5EtnYW9fw8
FjiDp+FEL0BxtI/gb5Nlg9DyvXeA7/eWJxNyPyV3ztfNgckTGQ7ZhCvBvjVb1BXS
LLkCE0JdR7L/bOWrz6f3qfp6xSuDWfmZ3rYTo2NFwbE9hvvwuRBEzSlMcy/ympyw
x87DXJdZNI7u+f0Y76Zoj/twmspRnm92vIEqgWm1JW/0M7uwN+8tyN8MuTxb9/bk
bx2O8uepiQCToi0AtSzZqpMvkV3kbnty5HN5jY1xaBVu7Ejy3/ew1Z1ZCkcgSUEl
sGrj6lWoNqdmKlCR0OhDhJB5sXGNy7nPD5gkvAATugNvVziLlTAso/kBEAg4WW6h
1ALkvd803mHSwCYw89jcXW27Dj/oje4t5OtK9U4NvA4ZgAl0+bqDyQ9aU+dGpNjv
miwvy90gkbcMBNiI1rOLns9WkMKTniBO4czSjwhQy+38uV6VqK0+NYhWteCC/P8g
cIv47K37dgih1s3O2z1/lGeSmZo4D1JlY+3YGRBu8Hzi46BFrajSjRROaBfCQPih
2UB9QJK3Pv9ZJaEmNMuQJkxMZGSMM6CMfCGbS0+sk10t8BhbTlTJk/tnaqxE6Zkv
s1Rwdc+vLfmetqmnvrjGhi+iEZfQc9coP+8qstfAQNFnU9aLukIyUZpUwSL8A38n
mR9wylDaQUu1lLaJIRyKxqKHR2GzsWhfAeog1xA9yLVRBycSaUhBfZ6Z38BWfAzh
Pac8ueOqnewcM+MzLSkrtNvU9Grpjpjb59cL63Gwz16YkCJSeijJwruy00PuXICq
46z+pzVzabx70MYugOILuDmLdT+fiwHVAKw9Alm7GM9vyaE+DfYZFAjQCdpakyuu
2lnCh0FVf1vfG5xMvPLjS6nVSI2/IQe/1YBiFr1KmtLUwuroiaclq6PfiTqrZ2KG
0ocL1vS07YzSmxX2928e62PoHKozsgd5gldqFAVx3nHu0tgDDTugu0lqeoQIYwAi
Uzk8sBceymlYztEzuAEtel//yoYHdjLlW7b4kyFY/cDSMSQpVcLfQe6RuJEaywRi
iNAxc2SRXsfkVAxmiaOVE/j7kHCAVice3wP8x0dEe1jL3Ir8HcoYcSS1NsxQRHK5
Fygq7ryNiKEMaFSqhqYyufSf2/Pwl47elPHpmx0QI6qo8JKpX22kKbH/NMs+yRjq
rPUMO9TpNzN+ckAN8ph0xWKhvx7rvZyVXf0xshfjjPIhKEDtmIyuJ6yFuRFmtBbT
47Ri7+C8j3akWF8WxFEcN81Qydu3IISGfd29OHnVMt7UY0/12Uyvn1JqJ/QYCh8D
Lu4eLdVcRdU+uHEak5ajnpsIXfkOHOvolCNyBFBmYQWAF1bnGD2YGv6lUqk6grWN
1o8XoRK1I2rE59gRijk1GhiTVekn50vhwL4AgbOJrk4PURMZKycpyPO3u2gzK7X3
ShcCJG3QxZjP2PbPH5YKbmt9aGYrnkSpWGkKpl/gMMYjQBRQwEfZAEOeoSnzsiv2
dsiSXXtQYU2woy4QuW5s9inUiv8EXpv6+cb1wXj6Jzo6FoUophJ48ZRhP+O/W22O
CUK7trT4IB1BKANRJ6B8FPad89xliTUPcS3JXF5ETJan732tDcYwQQMJ6/IyPaRQ
Hsgr/w6TA1X36CWZHLMGIQDOavyLRS7OwnAX7rvVmLe1Td3b8cJpJ2eDaJ4tqbF8
sYlDg9W139LnFpLcuQBDF/gNYhKaxB52dXsVz39IFSGarGnYiTObipI5RpJ/lqeO
nkJphcdYy51BvDgLuw3DR9gpd/YeqC8J+7RjK/0w5WuDRSy8RTeNmckKgAGI31Zp
GTTRUudkBj+3a3vvSe/0Qkh9KWMNKZ7MBFDk/8z/sHwXfqYwZ0kudmxMLjasWid8
YUqUeblA9sAGFdk+hg7IIhvpaVjFEJQXTcHbD+oWB4rkpD4xDGW3CfxdZKd4KlPd
1A6Gok89DFsQmYsT/w08QJ4FQSM8Ww02vrukOXcEFCwe+0dbmDKFXO8UwVaE7mEb
eJP0s9fv+FIHXJPhAD/FftugcHepaViW0HxBvYdwCl2euyg/Aa8LNZNZZHz4gb8V
8hRXqRSOXZPas5NEcy4wOyIMg6QDZ4ZL3mQPysIlPFDDoiSfIVfYYMPffCoZ/gfv
fk9X0gABhE4MrYcC3UPY5IJr2H/lF9wVRSWg33WEm7Kb7sovlIqn9e9NYkaKZ+ad
usSy+OP+IwG9O7kyd3IPxnrxcvHIbSvOYR4ajQZWsOUkMq8Yx5jyPHqc+VU9B76A
NK5Mh/U6AAktNVaFVaBvCBGccGPSMJ3qrmDGoAVcc0JUwji7Sfm+NaZIeTiOi08V
G5MiXX/r6f2w0DB9cxjzeEEQj5Gdu0lJ+5CFAu95Ao94jUdRy7yUzYk02oUMoaOy
FQ+UGPTlyCkMLETyB1ZfHYVaZZ7kxXmQazbEmg+OUu54k27FggJV8g7+cG6Gb78I
8nRVJtJAwv+2noO5W4jf+wGClkVjViIwpoZsYAaiw1kqdUq3LJnlK4QtMic4xy+G
hBhpBf+blbbxPmXCbiFZsw37vGloKygp2cb8K7lAIPlHt4aPt6w5CGoAPAY7wUAY
wgrFQ8dtjnAms8SQdET90kkU1DXVFsFi9fA/LTwcQ2eEOWWHzG2gzPRckajM3sF6
EYvbqldB6akyVsIvOWFE9llwlKlDOmCW7nk98nHcy2mFZ4QveNaEMXRPvhHwFY4G
1Rg1Mxzb0vfUrDo/2bj+e9z6l/EUt6HTatae/qui6i9DrCay2u8gaqu+pa+uxWxT
bJaKGFzFSmM+qXIk78GgZu+OjBtw6ZI0Y0w6nrdIXvC1H5etoj4DpY97smPK2AbB
ROrya6zCoVb1AZfQWwX7/dryKnTcpWnUjT2tyv2JZlVz9Uof2UXdx7J4Fyhq0zzo
iTyOu7b3wpd4jfai8eYyZyraj5fvR7K7FHPMxCv4hgQFON2ug4BDVHPTzZp2lH9F
o1zokqFFtblslbwdoJ3NGY6oZSJq4evEIcBfTPnfQtNAEL7hpcPV/80T2q+37Khy
oVspQDZQVBcJhAyHEAOpDEU8GgTDKSMLAOpc5GOews1TVCEY//c4p9etupU0ZLjU
SLhctbj3tGCakiZv/2yrPT/IGlZDXuAi3f8hQY1O4/vOmlOg8DJzLaWilOZj9mhk
erFTnMqmwwyjzdMgutD5lss3rETCUKJVatd6vbeN8ThlUwOwmt9/ZPacBBsJnkkI
LaivvmuHIvI0rJTl3aOG3jRmkpBP0vEERRwkipKbMkx9V812leyxnmLzwBvgjTvD
iiNeKyDiN2+HE+k8dr1O4FQA5bhqr+PHwgPUXWZv7t6UKU8jn4qE4APLc98srCWJ
sxIIe2Rf26llspX8FrpRBSPgn1HIaffh4jRGQxZWE93GKkrzVNRegk2LF9iCUqnP
IRn+en2jsyaLepwzHQUtXiMaNz2s536gKumcZAosfdAlJ6DdZFfQXKu3PV+gWDdZ
j+e2KwpvqAgNgelTuL0gGdqeaJhlyoEWAg99+Qy2EQcX9zV/FDjexEVhU7bcacTb
Qu/qNZToAikBEkMbHYIwhzE01rBzUCR21IXikq7M8JO9YEwOZLSqO+JFQo8QQO8x
2kvPwzQyai1nM9d/Jxk5jKQG8ZqHUKyE1IINwTyI0QC7US+cwnUQHmBBTlS5BI7t
hwXq92taM0WL/GVOJOIWBd2t5+8DnNniPa2f0jwGxK8fI/052coXksUcuQuQqG7B
IdwfPHXbTORxkGihK05MKpcp6qLyic7e82+MJXQL7EhcIBGI5aqE1IVYlNmGUGio
coqO1DhaR8JLKzzcEXqz8jwoIq4AG3tsCcWVfox4Y00xKUV6SbmFj3bD8m6C68t3
4MBrhBpjC5cD8fnTMGdhmnErKLyd9U3HrepYEo/7vwDl63gLad20mQEbo2oVfVMT
8XXk0+zuXnb6mXxv2h02UzXjGYjN2dJX6BcA8ffwqG8Ff2kiINxpNYj9QFJk6ic8
m6fqP5xiEmIPHsLiMwh5x6e6SjP/38kEuQ0zGpeO/C3KJ8e52S2hMAhqXlTcM+Fn
zkJb4jVMXNVdlHXZO4Jk4SHMgh+zUmTSY2vRUa3F0x+GIwOGHcZs62DNQic3Ypmm
QmEPDPBz+DzdUxlwZmCwsHjDJEU+WYwNEXrY1RCxtTssGGZR3WOQJjTqrFpAxZ5g
szoMSn7Nq8R5m18KMczAKSfH5dUS/CM7n+ddQ0WUl4Zoj5gv508Z+RtMC0q5QBaO
kmn84UbIeppNSvMyxWUjAVtJpxncCZzCZr6ttw+ccSxUxxE9zd+4P4GjtR7stfQF
0+Umc57Bn3HZpu5PLSBeRV/bu5yYJo4MBkJm1ef/wXzF72yjejaBiaPTs2lKAiJz
mfrdqbm75kBZ0CdRatfW37ZFJPiPeTAaVfLTmcWHVzSWVNaFJSVF6AMD/pvRaPN2
kBFWxMbzA1jqR8svAkVDyv2KEOqN1c3qGqKT5aahXUelyAh7dnBt+xIZZggiYvg1
OeknPrB2SloXzfDQgutIK3ERmz3AmFXxJpD/ivDaagZ0B3vUqwZias4wyprkjZdQ
RAsP2Aipuv/vcR5ftz81xnOYVUh5BKjzjF9+oKobGhCQwHA0iLHO4AwugQmar1bA
D15UjCKLCUL8v9KObJrwbFLcjFGUHo7swoLJBst7H1pm+oQia50KkWLpdj1R7KVb
yZhstMAMCxoe3chodF4DS0SQXRWNEf5MVCGWNWcXywGyCQ84r5r3GqWXNebWk1O8
eS76bU83RSaLrOoptGE8EBpexZhpB37hOc9YkzOOM9qEhyXGHYubMC712aN9Jbti
7TSXZv5Z4HbwU+oraqqSxR9vAOJL2ZVDg1DsVqkJhSr/pgISuFvK1I0vOIZbmn/2
9lgulQyqEBbYfENAR9qmi676ozvKXEHybh7j9fm89thbcmOd8AlKytW8mJGU6Nq/
KtRn/yla3D1A1KShrISQkYmaHwLIrmN/cvtOOHhPVbxoaOvFo6j1ny68IMK6CoSx
GX5jP6fpvLLAJXexJRRW0G2D3Czaw3KgpyXYHpwNgNzw9NenW7vGGhW+KMyyc+vZ
9TFaw6+uD1TedFuFJ4/qTTWlHVnmvu6zndkx2XsAMDZHZkFtDhCalFlFv6ulgoIf
58CRYPmuMVjPzG+QQqdmb1EoJCAUGBrm08UwNggtrZzPVdG2t7y5HwVwHmI9Vfyv
rYItexUdGcGAgGwCs34cWS/MnBY/KiewaGP84RuKJqJLOD0xth81BhVQtdWg4DNO
oMoxtdqEFLxus70TxqiE0oIcwoEtVJHu+QbaVUut6eAt26hzczSASJIz8uccalpv
5hYW8DJbvrozt81elXR5sms28OeRaS4UgZHu0dG7QP7UmTtHS4EERvR5+dTRUFXr
YYLORbqcv1r9pktozTG39x9JDauLRgHHvII3cYrGa0FQNtbQhntuJAj4BEy0Fams
kcdwOJIMBySc9nalwok9EWJ2E0F0UtEiajayfyBDQZ+Cw4hQvJ5IZDddRWRzrE0P
DbQVKL6a1S2gm7bXIfSFqb7StEokTSsZ38r3QRUbz1cTim0ySYqFrS1NiVcXLEsq
um5h8EqGxMvU4XUje43PTGajBPnwRKy4lqEudOP121/EvMC+CZ/Q0U4FxeN+e+oI
X8CeKPZo8aLpNXt272ItLvSfXXbLsjDGy58h0jE8t8pg0pC1xzAm1aJC9vLhgrsG
V36O4tkmRsbFQInO6DQ9mRtpD0Fs01qwLFKBMvmwu6EP/w7GboEY0huYKa8AR9E6
1Tt/LcSKMeRPISAbyyNAqNLv1Ie9Hgb980C2Q83256IYIErOCOv7q5c/D7cLc/UN
gLu6CyVDmEjFG+8x0T4dk83nPLPZtH0Cw+vB//np/4tXDhIJSklgEQs3e8u1a2xW
XdDWiWuQ1f6q/O45E4xsYhMj6c7VmUgROxny2nRCB0THxZ1nil7pLlnFIdfjA55u
BRMs3tWJyY9YpVyGQZd3f3M1Eb3BK93UOrTnUhc2m5PwkH4Gf9wnUgwh6YqdrwyL
79XJVuJ6km8JsA5h6HHAP9hKYD3AGy0ufZpdJ7SgTGGmTLxKvYQaJspt7ZwN15RN
kDNeUEQHB9jkc30AINdK4j77LTJGfxyHXIP1+4IGZXCYsKmPV2oRgoEgd6/u0kwD
FVdzs0IfZrFwFVq3saR2/obzG685eOzEODD0m6H1wrEqkHLE/7BbFiQeOqZnkmil
BL0vaVVvvN1T0v0/D7/QS2fe4A8dSGWWPyanAvY0CTu95wXAIkmyRVtmTKbj+AQn
VbEKCDTi2DJVpEzuaPW0bT3Edjpkh/PbsgzVIoV0CEiuXjBHGTcxb/3MWFeuAq4F
OpuKM2DyJeJgyGfy95YumNJHUaf9QCEkgL4SdjYtd+nzp9qEOANEYq+gQiQfFHd7
REyofx9D+ulglk1Hwq7fO4938SZoYQb1t4pCpLHKWcb9gETHNs13VDoj0LAfdkMG
h68kn5stcG8X5gkNZ2BrTDazs/scnvYiuEB8AI5H0HU18AvfVDQXVvSO0N51VeYl
SeNRsQbXGJT0G28j6X/RW+wZl07C3kUvLcsmKkiRx3eyGEP1fqXZM6XiMF625bMG
R4ZrQRiEf2zPwbW3WGTuj1EzY/tF33c1Vw+J5C0HZylCx9gD8imQW5J5ypYzxrgY
tgDWoPE+ABvHXxshWg6tICCNXqOLym7X2XceRG/BSnU0TS4u8pEc9aQLD9y1ZKbu
B0UfMCOtyJuYctGphIg8UBeo+/UAGcibxpkyIDvHX2NO5AAa0fquxBNTZZKE08Wz
a1MNlp2401Ynlu8Of3FC3EzKFuyMrDxNAjuvLai6Y9xNmEbvgFkTzpoHEwECDsbB
rReqnSeOcNZBK95UXc941TNT1dj1dwn/qBVXW9hWF1/Ckwj09pzASeRxEE2BhQZf
z/HD1iQSLho980Ch6ze3uBOj6W2GpVLB+IvFS9iSh6S1+TQfEB6gM/FxJQ+wucdy
aKLfUFHji6WQp35t5JRi2Tl/cA2pFZSFXQJTG0+zmTYsUV99SEyvkCWhdJndI6SC
lnPqh9BZBCXVLEXZ23bpKMXndMG37PBB6B+g1/s0opbMZW254oAAxPzxBlz6jDG9
I8oiZM9YlBz+izHGX7TyhvUaN7gBsfDxtvMszEWSHWQTpU8ErVHb5Vt4j5aPXxkr
L4HfR3V+6/O2GGCD3MeyDztY3UylNdFGsXs/rFM4eclF7OS+lZKQIvO7p3LsT+IH
lK56XKAuU3K4yn9dTfDa/berZ7lf9XF7ReBhAfFY2sx/mAZHtxFIAhOy9wReBj13
hS48UQ4L9DnZ1FrYpXmTSVEjCLtUctyiq5R2Wvr8Oco4a5jU1vGRWXoT926+1lEP
zDHZAygcWlkQM5bzLSl835B0NQQXnXKA7NWS8pvmUzhrPOenF4+qPGXwubRGGFzP
jT+U64aiQ7b7HKhFrG8XGdUSu+UJYrjUouX/FtqrCkNOaS2JkfEfaTLJZflKDqX9
LOmDIB0ooxE6qoWa9g+wjvZ2LmVupJpj27RY1VPaWbVRBrm9BVG0N5hOLVcM3r3N
wkZgvOoT94rdeces5khzAiWLuCBY2L740WeO1LIzQsO5eLpfpPBquFnv1TYhG3jE
cb6oQkSssS6aAaY5XhRoIrIePL7lnHqNkiRbMROAqB7fpulXTSpa9oha8BvO1q/5
vNUusxnaqjbxP8MaX5GQ95CnlATYETbLkZwL2q0x3rrHCCdWh9+Q8lzEEt4apx1P
SqDwe+M+tSDCr+zsHFqL8fgGUxIIap7pq2I6V8DwTksY09rD4YatZr7xj0ZpoeR4
7uSjtqis/HNugTJ/a8B/aHeiXCIMN4ATPFqtnFbntp2cZdAhKuh6IK7xzjBLFn4Y
JjgL5jEr04TjEvFmvyhIfSqbeXsBCwtm2eIZrGLhcVuEi6G4F+cvtER8EdG103AE
Kt1Q2JhzS6/Q2/vsbXG5tA6tUbVKE9mLThQLBbhzJqwjRYtLxC0yFXyaEZjqkXcr
xdgKHOSepQFN2MkuuM8ifxoZp3uaZLi8N4dmZl16p+C2LwPCPepOAQx5iiMJaT/i
cnQklhv9YfsCMqoJgdZo3kcwD7EAFYoY1YR9eobDb2oVdsHNkSBZ6IgAulLHdlT1
W8jZ7Hf+g9ahKJsttaWsyKDYiU2F5eMHVhBVMwkCNPcvWI++nuFDkNn6sBU0ZHiZ
q7k16vwQfqh8vn4Bf2KdZgu6pYzBlvVQjcC2yQTzmUvMbJi4CriXllBMT0QqddaR
khdg5mQCndw83TI6Szu2v+zk+bTNUreDk3w8ZzooAGqL9WZGv1KIWjs/3bWU5d44
0YSlZS7xMQT1BddJP4ZKIRR9DeuMim0SDtj4aRUuN32FiwniKtBtU0YlyTs/RRCa
cwfTIUvRnVpr1kyPC0SOH4/0IzpnzZu5BtgyXcZDlbAW3kA1/PnT7nMpT32gYINZ
V+C+JnAtap1aqOxllS/MaduKa3oDlBhQzkxT+lH+bJUAB7RH/U5/tmOsHwA9RIZS
Oxs5ucH936sPZ7jLdZojLvyzYsKU0g0zPYZnAITydmLNdEY+zsE/QAnNVh+//9k/
wkhghNUTVl77YxsZIi4ltKaYDw2pBLJkkmc46fV/YESznhnUxKsSmwXtmhZ9agjM
h6PvNdiPS+FKLPHgv4Rz7G00+k6gFBd6YAhFf3P0y0kkA1n3w0TY2xxVdX84T1j8
kC9eg8N+kGcm5BZze5NXRGWo9GrmWiUz2rcpSUgktetXObbSxq4uxZNzrdc/KYIQ
sxYzwt6uhUk+5AjoXyzdDyv6EHkE/4E7dW35E0bxfAJ/ggZrZWaBvQV/z8Q15Sct
yucsbGuVfeKVOcCqA0ue38IVYNXV27b/Vw/ASQb88zssV11vtzNeXR7gQUOt0Oxm
aOO/x0+OGCyHw+3o9TbeWGzMyPAkdy/jS/wyeunxWJbW77pO4nCEcsaY2dLJxr25
N6zpBY4lUlaBIPz9PqTnAsfwZtX9FPAArl/4KPbaucZj44YG/1HFmkDKgf+YvR+Z
X+jthzCx3F8RYeJjncg4htq/uuJsUjXAAZL1buzu28CzzPQe+StD6/9rBi/OO3td
sFaqW8OEYW4w6usi9V1wZTM1ae6h/gjMPL2UQ9nzAXdawGiy8mQ3ByRRMS8s6rBo
mduNvwK9VZlcCZemKHUXqBdn2KGFYgMvKRgC3nc092qhE+G2Xx60vdB5qIKD7oYh
1vsrzGv+X6De6x2tmQWO4eX+BfaqqvSnzL3a08jRkteiUAvBoXyX4V/so/QblP9v
EFkwmeCGtbzIA99hTEmHYFvlEpg80jp4vDklWqUCriRlZWlbXDgjSY38f+DsIWHI
sllLtsv1lc1o/lQiAdkL2sdVcI4LO6z8nbd939iTTbCIEn/PANBX2+PEFGMEgzsW
wOV76Idb3AW3/ZP9w2ZD8JU54scAn2FzBAJ5LRIGDD3C2E4ePmXPJHlzAO5fFf+C
OTfJzPXGmtp+vGHORy5UB4JXl3lz7Qag7++c3xqN/iR3UPVz0cYoK+KfrH7aCmye
nQagJ49r3879w/hnMm7SviOuprB3fhxSS20F2MRU0MfsyFjma3FkPJKpKiTUp/2U
yaGNfqjthOBtWaVJxiYXUP2KjXYvGklWFZMtnpOXaXEF+34oQ8e8Rf/DMFEj7nrj
plC3ZxTItIsouvOiCjXX38YjfpuBeQ32VeifEavq7c/QG3S0Z7NiwwWjZsuE9zqe
TgreqX0sGuJX+S4GNAMKXxnihZCHPEjXeuD8bakadgipRpMwV6K37x4WPTr2/NHu
IKpJUylvBdz3hUCr5AvvWZ/dx7JOZ8vZgae50KhUAUS+vrPEZsKHmw8lzlHAK5S1
yM2dapb6vkXJrgL1pZRv1nl1yeFPLsW7iZsyVTc8PcrbMA1E2EYD4SCsOhBXaPnO
7QAqRuKQHERg0k4BQwFwBT/hUENS9Z55SKz0aad04Sp1gi8bPbiBTVvM6ae7FdfP
BfQGHjGy0UreByBVxAcA3vRqnqXisdjeKcNpEA19qoNBLjw3q2zyrPUc5iWa+hYe
ui3E5Lch3vzMiHln+k17qGPG3gVGN/ZJlFzkYG4YRbVG+c1Z4JLZTV09CPzl4Mm3
lS/1KqXW93qf7oxy8OgqNMKEBpLeNfY8VKk/PcjyiIe3SCu8ZBpgezbRl1WCaqOL
FdGOjNmPO+tppXu47nx3QtzzPnoIFbDm4WUg7xoFINivAJzipjUTlK2iKOWi1Z4q
8ssppJATuZwMnOosnqXlI+WUUeQ6ImtqQqMU1XR8N0rmYX79FawbnCKJToJSwR3U
s3JjF3tTlyW1D5AAn9ktEgAsSR+YnZoEBJ+DBWbwJrPuFzKMDJTUESOVD1MYhS4n
aBFsap7yqu3nVUY1oLMdoXBTVVxMR6ir4GbBcD0aDMFzyII3aY3Hn3Q/5xoNMwo7
/y0ErjqmdbmIIGxA13hVFsGuFEGD/HjffChH2iLubp+THSZVA+OeiCQ+uGHEGkgU
QbDCkoPmowMaIK6DM995oRs1cCJ4ANATdXAyllTinQcVf1o8vtlq3+9LCtvooRib
CQvWPfd4VqYWX/MO6EeV9gcK8uTYvSG+2MKUMJ4wSI5gcn6klnuyxQ1QS6ihxUyi
rvi2x2c9ZpB107/eHHJjfK/usP3eXEf5VwCV3zz1EQEmVKU+3SDsKypVGuHdoANp
VaEjl2iXNtujIR1FkuWG/yPzdQz4XlSDMyLdmkl8XbGm1BbDEhex6aG5rfbrmOsO
tYHAOGnOOfzoKftHRRjOCBADdq9/oT3zk9ajllJbHaWqzs7IwPs4DgPWly45jJU1
UjeW5C8jJtmV+yar/+nxPhoMXaMDuvi+W0K8oDcpU9LuRHdy9XDHYmX7gOLXmZYn
n0TPFDuuUQ9FoSalo09w9/2GFZDgcN/9jmUT0XnLe0iEP4HCeWz+kSf6rnUy3ko7
8Fe2eSi7aY1Fpfvtq9daOUk+bPXoYdmDd+s9nBddoqfDC3gKQH72T4ufXM7U6hp9
79Pfd0XeG2LUBUiyiEVHF91m0OlOg3ooGQmN0Mzc3gA46j6WDWrLKK6qwftrHRR7
VcctHL6X/HzaonOsi+L/sYmerLyaCdgwzJcf6DWMiRS3x7scLCkVmV4QiepRbrjL
YkI/NunsdTYYVK/bUmxbFkSNN0q5T8fh3HpNZFLaffllcUZXXmZLTtuU3dLrV/Mm
vwNqy30KzfRUOfeHBOlHYe2Pb20x6mZmniqLI96vaSM/cJlMO4ufutyn+TpEZB5o
JV3IH61qlD9CmzjzJRH5RHP/pHDYVxC2GNm7Yz1ApBRMSmwddxHVbgsXo7urbDvY
SIrKoTbTPRZKHWLJWuiC7OAW6C1qlj2VizU9G7mbuOj7ZoZI/kEH9aepJJMKX70i
pktkHQKOdpfZefaLtFmX6FDloWfAdcTnTi1q7l543bB5rHa9BkcuthumDJHy0nnP
fQRHHVyZ9jl/UPQ6mv0xhzRv6m5xW4rbpKkPfzSoVZ+F69o6Alaxy80cZnmgW+/V
oPXYGTMK9dimA9L4blGCuCGsq90Lm6OjIAD0adxGc6WzTmuwOB7pjFzHYPOGQfLM
ukPM84Cl93t+awt4Jj3/dBHVs4EkN+N7gA0frNvJ7JUCKrjhHUtk2pYAhUZoR8F+
Lv9cqWYIqFSRlqUtdPuFFdKSKSMHZQUbqPlpjezf8wyB6Jq2FgGrt3pQaDUd5OVp
w9hiU1os8sBsmDPHs9eSnKEMlV409A2+6z0Mf8pM7m1rR7+trlqPHbW2ch7c2oLc
w7Tg87QW+zsLpl+1C5jX73jvgPgs1bwFAxlJUKIyavirSt0ifpTmrZ58T7KhP6MZ
oF2c123lScMymeAgXP/wKC7UcjlxWf2efS85EUPH1PlinQGWUm4gZnABOmLshIfV
qRKNpGaRMtQ3LIgsPpqg8XathynH8Bw4UUy9/jDOUshWjrefm9A2KPgkCND2g1a5
ajzh47rKzWVIPC0459+YqzBE+u3IkyNgAGooWBonBWhQAXzwFPjmieR+RUZo3PYf
wYEU6D8tH5ViejmcXujQ5Pos5CJH4xPcmzGZYsLTOLeauJMAML8ox1AUczmjBx3p
HedPM2vvcTxR/+CQn/tk0ZC72LCRLXPoeGdlAyORUiV3spagoWoBapuF79RnVLyW
cS5Ab8Y0gbv7QkW02SYSqo9u/fpiXIKcVBI+WZMv41+f97c6MfGe3M8jKzG3BAfc
Qnq1S/CMZaR6AgpOcxACjk/dgk/Gh0JTbdVF4w5DwVybiqfU3uMEUNpykNDWbfiD
MDsTBsZtLfQuFUkE+WZ52I/z7hV037Gy3eMj+d9zMmpW/1iBl/t5MrNyYf/ljEpl
nwM5wDNEsxpJsjBaVFSbgOQvsmWkGnE8R/E7//XOWoYzNXNWH73Ciqz500Qlczyg
gZwN71rNntl+Tr44X3+zMoq8c2t520Gw4yg2BhdkqVphja5MfavdGsq9u82hLMsN
Xas48R3oCOxpKMLKumcEtgU6XcRTu71z7LlrdJ9zatGB7u9Y00sM0pnVpsJ50V2t
uMk4A3rZg31Wh+EuNT1+UIT4JWXfUTtznBqkh0NO4slxFlj7oh5O9/NfCGp3Qcaf
g4Mamj8Ik63pa4fETvEOBMcU0cL7LEyQFJpIRB0LpRolhgZO/00lZs8eANJhIaKV
qaVKaekqx1gFV8sx1X5OU6Mp6rOxFpDZ4MXmTyQ2rWptGjSKV1wlM1UskzKmpDaX
o3VSz+JgEGBH1FFrlWFZ+oaWeyFbgA/Sl1cv02QR4DZ+WBp4pOSXpoBiaSicnfT7
IjU5xTVQ6KDIzc+OBZf2I+LeUO6IJDQTRwF0w5oiaYL2wc6W087Utt/7JztNlzvR
cLkMAawsnC/FrVSpTGvIfMUYF604i4gf45MhwUi7nt6eMh5yc/QbdRRi18GmwdIm
D4ez3FEwNvPXvMWalh5NGB/qR3Q/EaKFLNIVu1s+r5EesKljvyTIH7rBLuNntkNj
ek315TGEqV5ZayzEBJZq1xnZFHoULX2G5Zpt035yzdDjoqQj73ZF0yYAChuUcaAD
vJtfAn6CPvMne+5SxKA/iqBjk+s4YYOqaTEUG39XFqInQbLjzvDarxTT9i7XZ+5c
sViyC+07CtvPDL0UMuFU8pWYFIU2X3VR17P9mpxNICT+3y0pv4/o03GaHvuNzKBa
PWdg+wVgbL5aCWE6o2gQYw==
`pragma protect end_protected
