// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b7Bb2s8EM8jcOSvFZJdzNBeyR26YAmo/639ZCt9x+vzHGe3ly5TxHk6bh+UB0eQz
ADFJqvXSibgbgaoxnCvu6PJS/k5l/xiSKi8YJ4RHB1F+VvBCjdZlrm8k53rzMgwt
W0QDC0eevglMWG9p8jCKdmKQ/5k3T6T5Pplg/+bKfnA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10128)
bhCjiNgm/osWTNBIn6tgt45VqtFYEW+q2NDUEIUDywFnsVTDRxNFsw9RxpCF6I7D
vWnw+n8fLqc3xhO4VY6eZZD2HJkQGIasu4ExnSKBkUC7IDQRZ9rpTCfMLiTMCaOX
ZTmnu/dWhTbFhYUN6XMGH8/rfYvkMbt33xmgPJeAegxxRITVITjQDpphOoY9b5IL
OEeNAS1gNBQRsyl2qvZlC4OypT53dxOjouFPBtqLwPmiwtiNPlmbWyKyfR3BrGm7
ARcdWgTo9Ryi9oCgP6Su6TycKDRxfp75wDZ7uuOUAY/8HUmzwqjKtKKn9foPjHW/
1EtIjYs2UvN/eFI6l2SVD3PJe5GCJtJrC8Rxa/xXUhIZXQoTpW31MZv0IYC+OHTc
WJbw6XNhYO2R2H003OZ2pgxcTJhLLqmNyx321fYNmyyOK+TwHG695ikKyBoThoIY
fiY4pbCXVGXui1aqejjyIG+wMj8wjwF1Hh26QInC4XOgubVYe+8rsm7+PzMAImaH
t2HtJ2DtrkI4BajVPqeie4os4A8HVBTNGd7j4alMr0L5p6QZ8XOSFAFj2qZie2ks
H0XGpAgAILcqCl/I0RIQepjdaZgkxkPKlYCneYB1vyYOcevn3RBvg7xQNZZyMRTN
G0OCtxZ9cTkT4xeZP5cqmIxBq2EGx8qtEw4fdCxWjUZCgamfeoiDGwDk79muaMHR
M7ivB5tKwKTzheutZl88YlTFaYptNYsHp/Pnx/XBLa6aeNWHstfecgMyyqI2O6/u
wDzSjvxk2mszZOofEIXT2zPtsA1tnFzhTaQMxay+t55qiWkMgIBwhpR7RtdkBeTI
El3wtdw1ztOHZE1BampUew+nu5JInoYcdMPiKmRBbva8ULMg8wXVt7N/rDAgLDDm
pnHfmCHn4gRD3+5aQQlP4OAJeUfHVMxbPPvgjaRiTkrq2QkQ7Bpqt6MZR4oTGfuz
QKBQZ7gzEe5kjhHJq5EW5Z3bHlOaGUJWmjo9KTAQj7jgU424OOXHOUzWz1ZTnXTv
wDx60fYjEiG9LUbibciN/6ZiJSYUKAYjRzAjOf9Ilav5SFq8KmmTnvin7RGp44Tx
yd+5PREWR5ineheYhlNTj/hImQlgfNLoJN21g9/rDbArMROelmYubvv/M7PVxIs1
OFEjXv+Q8Io3lqb0zhTxzh7cM3BVJBU1+xV5JEXSxigsG3oBU+voI36PpWiPid7v
/LiYVOtfqLilubKGgqEBNFfz8+bP9hY8RNWJEz59rs0Akfo2KRHyVZ7icBdvuGv5
bFDUjPzb9v9AkEGQdnY7FKiQxDtVjkhSlF2wKgXbH3uamWmv1r3acm/mENy6cIF9
4gNMf+EsJCDShfDUvFQ2cJ8g+LPxcbrzXDmRMkfDF0kuVeUVyi+/dVHcO1iEWGOD
dzkWsY3IVP99XmLlIvRPn2mJuma39JGUqend1yc5HoP8Xjhg+iVhiMhQR63EAzv3
h9E1pLSHVRZKavqXmUnqrq35gKY/5JxNsRSDs+ocZ6J6kah2P2mtNX5GGA61QwyN
ftnTpfsH9OkcAj8bFwJR/hWctPeywFO2H3l3m2tM9WxlEaSps+X4XKCU9fzeTCGX
r/u0+2bDnOEj8SJHDF8CUt21XIAPm6A8aj/+rCMiPsUESel86YDW7wHRccbL7J7P
kLLQ2KCjyd1WcL5ZW1XP6BdCJAYlRfpMIP4JSPaKR9AioW9sl6OXgyWvgvr4Ycjv
4wJTS+lppcgYPmlRv186K+4I1PL9aumStF9hjmQlZQNgDRhgN3uM+Stlrket+MMb
uT1secydxdOhWtkLCe+nF/Mc0kYnCrMMGSF1eMo+WE2Nb33mvITxuTTxA52FDyxt
+cfcR1sXqRbjhF9tRkKkXMAqGCHLzRVQ17SVgnyB2PmVst4o0MXFOlR7/obCGtgi
7J6CdgatGiXjzb4VAERaMMgKfdAbLCjnACINiG7xu9ho+smWI10I1oS3HXgD86JP
EWo2Mu07hEF0ZKzrW3EvcVuKUt0ol79UARDmsILsj/mBaJE0ldDRwmPqzi0ENswo
vfyM34mJqip03OCGu5Q/RPLlfL5yWSWR/plj6sJCGi61z4REdi0nHR4oZ9teZVbu
1vJhwCjbhOy0imrZbNOD+kEuJ860HBYwXhthLFP2LFw6N/nsKCdGIGRcskLmTZ9M
/gikLtYGOGbrrpGdBJ8BwbL7j9ncPv7qlLRowumO9Dkt3TaFLW8ds3ASgxy6mcg0
JRGkOw9BR8aEhR57GS9tdQEfU5qWsuX136RQ3IasQpFX60nai4nx507+ZTssR3R1
zGVq8r+olKZHbTRTFC//m31mt+pNEX2ri5GL7rc3RvmZpWv30JIk5Dxy71GNqgx3
rV/Wx9soro4on6scClnG0d1CpsVqD9Ex6ga6nTRQ4wa0gIg0c86rhII6PcRKtUmx
bj5zIbcHmXk9mCr71ezpPM9Kfbjw4Y+ArUkfCuubPoGmldx1ghm9G5007Aun3bvB
Ru3dPiblRqX9tX3lX7GOIAEmgAlpk6BNuNW9MNyPbZBqLDdVRvHNh4PdoHzhWG41
rtUChjhKY5XtI+bVBzOMWtgwEIZrh5r7NKMKjQNA3YzfDvWFQshnjLPSyUR7fZ9F
VCmTv3V1g9uTxPhKlWx7/qF+Hgz65dW9u9sHIA6us96Q7eabP0c2cqHgMeFMAlfd
WgOzI8YTw5XWGkRfIGsUUu6c7KQ786sycUYfY8AUpJdbcDOovBxms/64T/5hVALu
wOK7Rb7B+IGNV7tm0Z8LjaMm44jNgCgJdqIf6A/icoOB0eheK66Zg2Wgm+/JA4jx
OKvp3qt1BfrdWopslvbiJUcmhVnvX73RXqCda/fCJ4VVp45KHzW9Sk4qaIvrM9qD
ERI99WP01DP5hJ4WW/TSSCWDSR69Cbu2OhGsN7Dc3KcBM6NgZeMC1gYWmOoDG+ss
7rtmi8W4VZwwpXfXnvZdgrR1Ib3YvbPHKYKbCGiLjhFQPPzeNkL0lcxqQ/GBijMW
WUwLqGd4Jv2bxKkF3BMA6waC6b/joe9zxlNtw33dx0KLWJ6DzOP38rOpIQf5+wOD
wUV8Aw/JcWcjFWWnZHoLKgWtSJX8megClPJhUhqN575+8cmjIVdyaDgabhyGoVu/
skvT9F2ryqMRMuoKdBsmLm0wuf8Erupmsx0+4IpM6cFruBStXPVSDsgh7AVKdCtY
HFRFvZCM6kpLNUEvEUYT0nShdVv6EFnwZ+/dHGrNJr9yTqKMl0+u6E/NuLNcULtj
rmanHHM30qgk+6ex+dEFITdoHhSVR81dA0Ja49zEXu4ZhzyFSnVCaEkrVagSjpMD
PKx0gdtZAtTk5ckTSxyQCrd5CvbEMrZfkXkEg6oH0xWNu/2uvAxliBOmO5KNmCvK
Ie1BU223g9oe8nUUDEI4+Qcr8pSuG4YLNDK6f7iK4bE2fyM1QHw3wz/EYnMXE5iT
/1lxP0D+RVnSWAwFsCHpDE5TYjZs4ENRtqxRobN2V+DJrLAAEiy5IE8noDZWQtWC
R49nixd51eaorzGsxEWJrmufYMXiKAyyNVrFhEY7ItsQPfO37jqRcsPepgbW/oHz
KwZZWa4NEJUng7X1vOySNqsi4E3vnd83AoFlKMEY1NZfpAQjU8hkZpeBghHifuMv
dCc+YZKg2vEDImIkZnhWLqJrjoiD+omhTsAR6zFB6Y1utN/euFm9kX1SxmZimzzu
Gy6J5yt4rXuoTl03u1wc2c8+GSpJsnOpUeYJ+f/JnMJmRcXxkgcij8liTezuz64W
VLua4CTtrDErw5mXSgTcEVSCxN2mWAmkgomGR2j8mqqMMFMw/5W8JdMw9qU0hf4G
nYbFA/zOfleZhjAqDKBm1VdEQ8MEZwXEJzsPz/hpqHs7D3FVJRtElUwCNhI9w0fO
IUhRkKk086vEWogiCeg6wefjlbpZiLzP07HaUcu6lLC1oYmRfSoKPsbhCybJaoZo
LSYhUgxXAtODuUQ8fBYFi2b5G0xhNbpM7uF4ae3WravaAD/ywDgXgfS4jv1dxOf0
mkx+ikmHdL1SyrU81RW6SIRf7/3QxDI23oyTGv8taRJ7+DANdr1X0DgQAB1ORw0O
P+UmfIGsmrwy7MlSxWwgU4FfvOHXr0EM2wtBQxGPOEiDQxSG6p8CbN4+148GcNvB
+mJz66s7cO/rVQ9+RgPsrmVfQi9Dpyke3v8LqLXwHS1r3CEgAUCd6tKaHWTvi0KU
tnP82XsZEp9uRD3Wk0613YcEjRJ4hz/Suj6VYX/DfE9l30srgrirC7KCyoctdFl0
l6HUbKfA6Otu/CARNdU87dIk2QFOVbf91pp0mXSpspQvqbYv++Gddmk0a81ZNYsH
+nVmJLWCIL/W221arLyUvp+kdMb4IRZZWWVjJpjNRrVGhyNgHnpbdr9fmGA84BY/
V8083mTL9krl6jIhNmm4js4s73triiQXice3d6qMfZ/0ZdXsSG48f9GdpUy2o89x
r5RWG1mt94Dx7g06kZXdrFVXpeKznpmIR558z/eMf5GNZCoSU3BuYPf9Gu1c2Nnj
abNCFAD0gIWw7s5Jjfp6oaFm0RQ3TUwX/qwK69vn7dNadTZGbMKvW+PpwqqA0bhF
57HDe1zO+oXuWMFAC7yGLEuLShtn7t6s+eZ3Le5iXKhttwOglVZsXJSWUQWqwNpe
kJ4ZhxmwRoHLe6zQ8nAfIG4Dji3CFE0BqaYT7FTHGV7PR++VQaa7rIkwKkZYTG1E
lj0inHE3+L4Z2LXEFjJ8QnviOxzuYYmDk7Zz47yPG/7AeFI2KSHyZBgFOGeXCGWz
FZ0x/b6H4S6kOltpuMrSvK7MiE/z5ScZfnpJJZM5AWfvvNaNeY+6hG7iiNPR8MzF
mQyGvvWcPv6DGSaHCY7rAnWTLJq63U+3dHyjuOyrYD7Ionamii68jSkz9a4Zz4Td
q+PmU9vq3MxFaT+ckAt9dEtt9UwxR+6L6OGEdbiBMB0xY/KaG180DDaszAbT7CSS
17DukiNhLnuWPMJaJa/5pkkveUMQhq/PJ4aCt2sUmNTtaQ84xZCT2P1tS/Ejz/Rp
Rr4OQsJYx33te7ZhWSuTnQD6bW685FLC68JLCXsAH8NiRoq/Ux2fYVXF1J2F4KzM
0xr3F+LTYnJnhqko4OwTES7ASgZVsszQHwAvKLfCyFuRu6YLd+dvHBgxjFOEhdC8
yj0/JjTDQPalFVLWIh5mSds6lDRYsQiYR820JEW7niIy7sl+YBXR86cGEjWVpLiR
vY/iIZm5xX0J+SYWJ0/I+pFZco4WEWESuquDlYGdwEA8GtDfLSI0IR3/0aaQ6/EO
WSisKmylaWFXysnGAgDDQYTEqy5jj32dHrx0No+fCeftcUK3Hnyb4x8CbkYNreET
ihon6jApv9AHrBTlIuQDwZMQSLPsa4bdWd2hxi5g8RsV0Wqtz/WJDfdV4+h3IuSs
rg4emT5gkxImT1zd51ZAlVFg7GwfFR78UWbCfX6rjY6ASq1lPXhwA34P9qloyyJ3
aeG7pgS4IgYTrmUKj8ULh1OPJOB3krp9ZGLZDDPJFA0joV08BQbsTjIW/h86hInf
bAaEYOJuGNfuGJFHZqLBhm92OKvwK1mTFDvSwggkWDn1DYQoBXn8whhO7lKB55W5
lxJJjPg6yEoGjt6Aw/a9JXgeX+7XyylPARS43QyDP8H9p/AoGyjeoDBgjEykV4yM
3mCjcu05U0HBxjf9pMAPdyR1Eu3rRLYQ2tx7SLmgrQ7CWemKJ/9gliaXz4hozwKj
OLSSlcYjiVLUSd/MhCqQEffknvE5MC0GWW/zx8+Rbab/iBLGqusbojRk8ve/Haw8
Tk/JCGe/Dzg4EpGJWUVaVLFIsFK7tLF4HabW1MSqobqN8bPBw1G4alzm7xQVQxe6
zJdWmJ9Im1cpddbaTGWah40WYrFvHccwt0cSV4CSQTsXA5OAw0ZGh+4ZEfMC/7Bc
LUSX3ZRDgM4FcL/+cZOTsH0Ix6WSEOEv7gDBFg0EIdhRXZ5Z8S33cf/2DTDegsFT
I9kROdpyiRkCek63m3R9XM41Wv2hJwlqjJYo95s2OB7olN01aieqt9hp2fJauCWt
/Fm5KBxUAkcFJf1o4uT54ebfatK6xCTA+MF835o4s4GUIC+Il30jTpwBWL8bDujG
LncC6lMWc1CeHd60X2I4aBs75Xe+fCI9P8ib7Cjf06K3WbyXNG8PJ1EK5wPsgG28
ImF1rZLEm9IOxq0JRdRtYK9W/pxtzIu//Sw4AER++tm1DNTm3D6Swx7Cl+/b0GkW
S4M/LWG3X5y71V891cQHa+c/fTAD/fbL1c7+8LdZKZHOoQp6WszFAWegYHyi74iw
ZXPKTVK8opndzJUAYLZ57tvGMrlnyW5o5GpvAmzSmN5C1i7NImqaV+Co/wny32zE
+vxgZZfgqysE6FL2Dk1ssGSDW1YipNrCPJn7vK3jAbMyjRP4XDKWp9uT8SWJ4LnD
gAicI+4dltNGa8mxTT5r1iEFg3yb54yZ94nG9Rca1vi851U9dv93bah7YdZ83K7S
6AoiU/zITelqvkIF1AZQZcxJKvGgXigmQR4U0xZDdQdGYGu3wsnjm7KgTTmbXsJY
MTqcWvtimOMzKj52FcUmMNep9b1W/aOB4e0tgtqHmuR44Yg5WOPRh8npV9Gar8/9
wLO9VWx4htxVI2hAFaKSQDSfyvFpXbnQkzz9DLOKTV9RkMd8LYpcdAtInR7sjjXq
c1B7fmpg2mA/m3YbQrLci+jAvDuDe/ldWXcUfag6TsYbbknL/2Z2t8g6Rl2/1S0I
looEXvdtz04sxCXm3K2nXVEoUkT9f8HKS3aHpLVsy3SE6HKcl09pdviFvKtL2Jee
sfMoWSnk1a7HkrGdiAQEkBhmqqjxswhQ91mQLOUtv+osVHRts9bnEpvBnv15SZgW
vDWSNOUcaEw/iDts05CmjbNHsS/dDDhdbiVB0JokEA7kYnm7Iru8JOdMfvjhzeuO
AdUAggzDhtEcXPsNkeg/aJWY1Row6ZyFk1arAUe3eVYvdXxu+/7Tyu9D/ybdESTt
cHCc3gD5tDcjGSUe2TnzYHLf+2xhOJNoExKSICWFVJ+P+Ypn0n7vwqpdP9F5+TVL
0V97deN8fbniugP5TPYPhQOOlP6vE+aAIJqVyUxJnE9e444QR3sY6uH5f/DsERss
+Ku/77JUvsUKEP2dKWJ5ocK7kWAwiIJD2n7AUAuC7ReuImPGrgb4biVkIzdIgKGm
fnKLIXg9E0FgPqOfqQrCm12KZTnp4D3Nh64VurDZ8+lxZCbkq+OKsuHJ3K46vTXR
4fCab8UtLIs1XBtg72xSpgCzYxltBb8di8Nsu+5m12lS3Uuw9eks7MTiZvKnz4Cs
h3l5jh/BSIAD1A8j4B9cCr8+qRpJTnRlB/TAqy59g3M3Q+Em5rRpGv2DRqm3jgKZ
E1ghWLvBKnPN9f4j0/i7PAHJ4/cwjTKLBhaF03hr6VJs+l6EYyR6oHA5QCOZNlzh
I2X3zw2h3+UAULzqY268Y15Cw/D7Payi0k+R2QEDGSLlPo+n5/VQ/1KFV9V7U1Zb
R7T3mhzCv5DMPyi4LWTtie1BH+MlT8s4EOIouwtUKmfJVV3ajR3qkAcdjFZYdzJG
DodIObjK8yVGhVrc6iBdshAP1uHtceIL4ra+qXzDojPs3eH+Jd/WoLt3e5vPtKh7
/TmLGGC6V3OzcmvXK6UURsdQmwc9j8gghKhRrh32vOXgngF6WovmKQUs2NIz85GY
U8YQXKVzWbxzhHsTK176qsRIKHQKbow5V31Q7OJ1k3cooPb21Z5IHQp/wtWuKSbX
s8/ZVkkEwT4SamJYRxQmBXHxH027bSnUH4mzMjL8IrSXHjG4sb5vvowAxtNiioa3
+j083JFJIoP8YSc1lTR9Len21dV84ZUHbhmio2EuWLxdNimzIT+uyYMMITcs8ZQ4
c8B/dhZxKKzQVXd3jRmy3JKohJAj8nEiDsd8o/8rqMq+NnjWD1Dj69Y9LdvzrEjH
JCMYgO50lhSuxILaxQdAvFxi+qsnQ/BHj8Mvfg+KNDsiiNhPIRxMZ3Pte4hFI6ZQ
BAMINA9+6nCD1o2HED3CEsDfxkArXeJWCmU3T5/y2Zaz9XbBogu96V/RAKK9C9DH
z25IkrhEZzCTiQC2UJsUu67/nXhYjkd9yo3JhirrIJ5S7QIHV7oI0KDXfXBlvcE+
bIRVr4TwCda5Lqg1ryolxOhcP+4f2MUFAvZRHfca57HFpEBcnYiEghNho0nI7kSC
Yx3c6sljd02VUyDEnktarAWowF+IJOB4nwCtMG0fIgcQ4tQ+RxFUoo00JjSQ000n
HP3SVbZVl0K2BojKipPdimzgExk62mC3Ag7po7PBEPhJQ8yH2SBKDndzd0HeRS2c
zcPI5AyD7eUrFjhBSX8HRzWlXTCiGk9AY+zWM1RjDNfKmHmgeMz1upBltpVcGlDi
2wfvGCUykyBOR+17oV69R3ur3sQR8IVwMWqcc8zpOQGMeDsXBJRsUCIvbccD+qkJ
0amAFav7w1Be1McvB2Ayq2HpF7qYW+4caajwVqPYJJJRo/r9fTfK6NmjjbqaimZk
w4+Cuh9R91mfcBuZtUzLWyteesTN3sanp17qbyex5wjPk8amfNd0aD5BcIkbK/KB
xo7Z79W23A3723Dmi1GMBMPCPydDy2gWGZ/lY2Q4wxzCtdIS1kZFQwwNwQpQE/2a
+9mNkaGOCKxdMqelezSqu1nKuY0nIswBrDjpalsMIlXoDaJ2lmQGgWmXbvF/EF7u
MGOTiVVOc94SCrkGv8n+++T3iYL14RtZI18CMh6FG3TtHvKi7T0mL9ogwte4IK0K
rn47LxQvzoURRhdk8ad931HfCHgu18Uf/A8Qs+GblXN79O3N/hirYqWNH3A9YC74
3YjCrE03S195vNUBubk5sLm37yT5HKmLB5NHezdf0bB4RFm5X+UHWrJ47HdRx4mx
GvOMIXzBzShvY/eMLeKQeGgZODDq+SO6VrjfmAMfhA+DMWpjb0AaeyoJgG6jy43I
gWSX3HWAFMN3KgYNw5lagNSxAlixqJXZkwZIZxB3LLA4hyIDOsXBmbFGQwLPHDLc
tAyEliaERObecVJCFoQGaLM4Gwgos6hpSZPNiOMllRx5nvuiOur05wBDZqB3JPgN
xLA6H3nr+EkshSCMG/YNLstnqNzzwTcdTwZWDUDcszyJCjRSl1/xKEPuDopyxqdL
LCFSVxbi+XHg4lQ4njZFEYDgoqi2eca10CIXj5igwt3XtMZiCuTWwABux20kOJB6
OGdnxcSNk0N9t8HkpNWXHbPgsoyfJb5qQ1G31vbQMCpcRBXkUqLa3He5meUQKE7P
tHqIxByUZHintGpsNVqvuJXFk4qvKK16egZfDEq18son6NH7aoJURXPPUxFkdAxW
0Ch3YABD4q7LXJroyrNx9uMycF/JEi0WGQwLTyW6D/TNN0EO+WYwGInTyYbBylg7
lwCtm5cN/aiqM87OVE36cw/1UNO2fpolOQK/+VMBM2uuIeB/fnYI5GnkQOv30zXN
+KZPtGnOatmr0pEc/sd7CtsbrXVZrsbHLDtxq4aZt+1i51wvk9+adbuMBMKdekMK
RD/w3xtTaJK4e0GpaolYkLIn6Xi1SfVo+SrmIbwg97LdghliQn1tegicbKCoMKr5
wpQ2RFFjWsMu7/wPdndVArMcuJI+2kCUAEc+Ofb7nJ59RNekbyHwNMyttdyT6OtS
cP/28rOlg4GoWvvCGsfK7ZCWq5qNL8x+xpJlkJJxxIXIAbBHgxMw8OeyFG9hNLdp
7cxjLgHIuhlQno0zdKJS4tKbWQdOfLUFwInAelB7+uDXMXeuCHEx96hej1cnftzD
JXyCkNEFVzqfRUmxRedRiN2Sa4pwK+6PC8fRrjqFeqlDaAZmw7DmhWOTluY1nHCv
EKycEQAZ2/EM1UllGuIVFQemm+oh1GitqlBmZTprrnCTkDuLj2AhHA1CXFdQT1Xy
2/ctdzpUkWAx/tpjICIbWR5Wse94d3O09vAbcIIV7PdSP4cOXzGQJ9PcFK3GhFLp
jnWsVMi6cxrU4osNXwxeUcU8XiJo0Hl6rL1S6+lWGuy5uKjTeyP8QiJ4Wf2ea/dt
fe7DfgmbA32w4ewNxpFnx9ufVaBAKWLErDiqdphtpaLwBKvVRW5S36N1yx3hHRdQ
d/99EMZE5aBQD0R8XgMv0sSUMC4np9MbLbgIuYdTjtQ/zGcEHZfABvnXZvzVJKQ6
BkVwRJeGPQP9LU1Dw5aoNtxy9GtRUOWh7HW99DFCf519cPu6TJfTe02fqnut+IUG
KIgjKt/5/puieiZpXDtOqJJxddpqMMobA48tXgJ1VT3aJ83O3XXINgUPzbOaCH1v
VXeQE70xn19Afgo4bmr9YdDZomcKB78UDo+ccPaz4JZdKRNdpQejR/rS7zZUvzid
5spH0Um1d3FCMYnlfIwXtzeosuX/wf89Ou91Wgxcnd5WUNYn2QCNG8nwHaUD2GPs
zUa/AzKnwM7KPA+6lpuQ0gpbwErmLbsm7hNlR3JK9hzFTkCfztmcluphv0/TyxLs
CZxIyyFSNgHKDUJA7/VqvgFdPnxoxwxF3jieQA9nPSWsKQjo4rjalaVoMNNsdBEk
BzncRZ2HnmB0xJ/Vil12EMZk6IGebzAQRCCsl/n3x/oalWTYQf0EeD4diCEO7vpT
4QfFWhCsB6Ot4irPLmVHr5OBJ7JXOZYvq7jNEneyV53t/vi5beV9IDOtkAG30TmV
RptVt6ng49eP5PZgqCg0E5UXQUMEL3B3lRJ9BvQeGil+zfpWepSPReH2kChdPGEH
TQtIKI/UKcKmBuBfovbWrc6EMTBU5YGWLAB453FZ/OvjwyKNmAsjqsl0kagmGA8e
syo75QOYQEe97o5OGwHlhC8u/onjnQ6ZNy8qdH+u/Hy4ST4dg3SoiKKScVjj2Y0w
eR47aB+sZTZ9VJvYg5QwjY58pLWlE9M1tI5PrEdl2oFOyJb3fhUT3DZb/KNnn9m8
iBrccQmsXYzvfUQHIWBrH/Ax9iqr0MaLlvOja2DfL6wDpOsGP9eBW4IdAzbJLI0+
AemNiH7e7tmDQr4tgqjKhXWkdptLNkTGxoOLwTpj5sUl4eYqGdVuB01FKsWm3/G6
nAKxGdp1y/NgLhtizOxGf0dWuz8ULxOauqlNIke3b2lq3WvHBlUy4Ga7C9vKB29Q
jGY2piz0uZ+dlgP2Cgibd69fcF3T/PrjwZVDB9Zje8VsqCM1lhqZY+j/ioDwq+GM
LDEgzHXmzgmFapN8qXsdJIf7Fwo6lAWmMZ4RC3TKSzbXvvGGiJbffZMd/ypebtZG
0PTuj7mjjjbLF/OV5W8aSSTyCMqFUXpI8iG2ydsZxbH8ff639GqD8kWH8vETGPUh
cvli6zHyZgwRkK01+l+5tsqAKbhbc5wBkN6cBkU98FaikAQk/b+4COBIKeJFQKeb
tmCVoIP/P9P3W0GMxdSvCjchkCfejpwFf2/S/Hivj2Sv3XX1WfRtyWtV19Qh6kqH
HxTJQNICKEQV1AvoGPnr3YDUy4HtQ0CWaknr8m0OK3dglemvIOmb0sL3Jqjx/N6h
lW4ZUbhHS1Yh+Zdk99h904bLRZ1eVCnZ8Xfy+xNBapnypsCRbTzQQS3Mj7r+1igq
M8md0lZijgNjpo2k7Lkm3zAKhsdZphnstAxipDXMi48RgG0sYaKr3VbpupCYVMGA
b+5S9hFwtgIeeIaBVfH4VvYo3JJJms6IuyYIO8Op40ylXG0vDtKCraH/6Y37A5JC
W/cZlNmciN8uuG/nS8bGYCsu0l6PsK/JOxZDSheZ4bals3cdAoOPZnPxUVJ/skOE
JczlbmG20y8UU9cQQ78NoLhh81UswMr1+Y9Ujc/nwwVON2io426K7nfWgL3ueWSO
YMueicMBvkAD1GtorGt6Kq7QrzVbiwMaX7N4UJUJznp1oEqrdCL08+xB4yk+Imj/
XnKD6hQaw9cNcjbrZj54zus1Yc9zGsynn22nNJKJDq+Y4dudM8Of2WFUnHDc3rsp
MTgoCTcxLilcR38YfiZ73bwQeZFj4S/f7GT09r0jsmqCzq/ONsL3F5i7GizcKu8y
5VpEGW5DfcEyEXqfrvOBR6JegQGyqbgGiJCj918yG5woyk04+i5IGF8L4SaT4w0n
ebEDMtGbUM1ox+M8nKd+8Ck2mq1Iv2w3d0DYJ0g8rD2s+izotXtuJ5o+h+ALptJ2
b+T19b/yyR45Ckp1ggas/a0F07v3ycay3y5YdF9L8sdccBUiJWN4Ld7YvBigLHsX
4O5Jl9mljJliKeKWa2HeGYACxP9tR2KtB2H6ynb7h6IxkMCY6kBXYl9WHEjslO20
rd8guSULINBb6SVaD3pZmsAtVTrjQ87vIN7ftkPcdHo21Hi/nMa+O93uqBIDlU87
IF+Oq+p8y5nHhzyDLRzz+eQnSzXGq5VTWy6z/fH0W3MlT5Ho0z5bcoe3ilCNNz4m
9c+bwLd1NteeWHLJgzsZXOUqUd643/cSDXAQSdx2VDB+Qp0RumMJnltr8JEPUwym
xn5ios8brQwZjnHlcPht/2DS9/InCqi5eukvcEFFouyQDkb56Gib8mHDTQbXzPdF
JCq7falhicpql/EZhKjf1A++ymYrFdCBom9w5QUoQ6CofsidQwJrIL63HYShELau
nDLn7F4kAWbRwbeGrOoNPt4XYbCvgOvilk18P2Vcdgm7Z+blJmwGqK70N37RMuqt
cqVkYCO35Nuwj8TvCqt6xZdGdcOrY7oF3MJe5WHbCvcAA2Ek1dqrNXJ7LwTXIogh
kNBe5F7ECPN8mo5fODvv6/05uVf7pEB1t8fg1FFarzYuRixuVNzPbTRKVvXZ9G1O
xIcRacCwLASUO7saS2pEVEr4Si+4u53J4flOPKGqWuQhtwfcXz+75Zon82/3kTjn
UvcntP9B9mE3L1m2RwgRRXUhi8f1Frd3Sqx4CbUSiGUmDmPjPUuHQsm87PK1+25b
IaegErRVLuALtA9m7bx3eCTvBfNQwJho+1qECay02OuUdV+rRqq72Bo+FccMLCm6
3MtZdMT6Ae7uPC8MoS6pt7y4awT92Hzb7IgaAFJvePbFJz0U3qXQxhJktMQy68o/
o4/GhVunSgxQXTiLrQhDLsgwxiOYToaLoOi/k909wxCREIdLp6EWezhZ2e8TAjeU
U8QSOSuknVPObNDndmOH72ZmC61x1ZNsGfzdxXO+9lPjCtGZsHSd5gXD0FKbei7h
xZTag1yjEL/DuXfTuSBtoCuThdvTYfw86rZYqkvKD9StEqAqvz9bvXdXP9SLDHxJ
lgA6hywA1MRKUWtZM62t+GctCaozpGY/QzchvhAGc1sWrAq1Vlfjl68HnPcQetJR
T4gZEUY45QZ8jmCMjg2LvoWvGiMS5P4Ogvudkgx4SKlzE3bFmfevxQKgPvbSWzoa
tCCJz6rkoodS9FXm0JMwK7DiXnLshmUmcT7KHmV0l9uFePndM39OFXOf+pjB6C1Z
`pragma protect end_protected
