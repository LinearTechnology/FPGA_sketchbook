// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TAYA6EG3dAc90heVGMvrA+JILLlC73NKFZt8XY7cGLGG1Eb6hAfoor7DXroK+ijW
6FIkmCae0u8zYAc2kTk2N1FxA8/61qiHxTv4uQLb4uH5lG7t2CsY0l+38ZMXDRG/
xxL/B7aydrl9Fb8dvWb2MZH7g/VW/3YTd3c2ZhJ8vr0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12304)
2XiiIAYJTASZoYJDEm4cJWPsTqQrc/RTHBNC0rvlEoVgUUMXCL0GgOsDcfLwo/3h
qYLbCaSK3AvxHJQOEJN8xJbUYC6lPSBXstb4cMUXZKg7/JCKogSW+zspUHmKHIVQ
yfyMVzI2Ipj74FdgBnlaKv6yub18JqD2ecC4Fwni+5P8SiA8FkiuDNjKDNpeG7vT
kUJABrePGNgH7ZnKwhV+XLc6AEZKrHEqEthnTkq31Sm6tj1R6YelW2OuTuqfZL45
RgaWXl21BijOyRlA4UVIkjiwwRPoBFAGuWboA1FjWKXwJUZ8yp2R1luY/6AffbET
UIdcqsQXOdBNR57FFp4Np0/h1ggrX2v4qErU0rFeHoW+h8PpquQJGACf4HlU/yKj
UAvXWeN5fq0lyKs1ZhQyN/+24IBI/dR7gXQQ4N6ACHavwBOf69tBtVSmn4LYsYJO
1PewU+rCTgEUIoezTuTtowBhlRKkCIuDRG/XRHI5wQjtM8Kt64sThVtaE1l84NkP
nKxIkFuOrNXGXhBUmqDEif7GmjT1CDbifPHt2eWbdThFNuQS8MGFDygMK5G9C1Ao
VjnB2YAe0ZzCxfcl1dDM6mZVEmBOd1LwK/RTBZB5IKbl4sDQvZay4G9Qmxg1vnrF
q3+pvdVkAX23SDaIElfd4JiXnV0kotBbUkitWt10Vol4tFFHIZCjEq6uVHZsp4bO
9zC6wC400b8wnCSJADi7Ea10s8KOJKefijVMPdj/wjuNWpwmNfl3fxbRXwZBrmwq
/wEzLoDv9eSzHhqe/YDv+suXSdJ6lqlcwD2ZKcSic+nGZO+CUW3y6koVtKrAfbdm
2Rc/kIhRcieiTWbpTFhqLlns9NkHLsBnmR0mVpiWn7cqm8dK87TsIK+RI2g08wsT
JJkp1tYG/7dGfSQCeUZ3G2ieyHGj7kPSYBAzx/G8HcVZM1CBDILT122pTC6Gwzdg
LsSJZnCyyIvWWGFuSO/5Yp3ikARqvDgAOMFLRiAviVPJT9tQwLknFEMjkRyXfGW5
FHbArBHQkDK98WW8A362HxtSTBd0oP/9BNeERz+Ivb3hWaGxtWOfd2ojDWMQJat7
iEQj6Ui9qomPmsDa+fbeeo9T+nGf13Kh+F8blqW8xU957AXchFo7tnD+bGvoLLqs
cYxpwg6nh74DQgvxbnkOY5yWvO1Y3uuPXGaH3croTHIKGI5H9ssT8YbK85KLmIwe
nK8PuzH2+kXPn8ZXewg90KlO5ypLK1PKaSB0KayvZ5FBxFimuT8fdoBWTktppUz1
yLVYgxrnlB551w+brclwHP+98ufzfOAPJ0/h0Lk9BaW88eLD7Bb69OTJ+N8IYvBd
JzGygZkdXOjEPRRZRpNM98pWN0ZoQNz7FAqcN3BWGqJ9mllifjFrhlhXxIERbc2j
KXhWVp7YdiLxbM+v0Z2x1d3qZfXr244va5G/ucqExYIIOQPQqmnDVVvQcDYQ/HBA
YmYy0TDSpp+QHH+3WixpBfpIKsRCQ/4dh3PSucpqKtFo7xRhSR16JivnfZzr4Dxl
Qv6V01oyleg6DZF1J4N3aaIMQKTq9n91RiAUaRs3VIiwFQrO+H9vkQgvF+BTyIO5
3BpU7RVRjw0Q3eUq6cMLGL4yad+tl7wmlHoczQgyi/eULt10O8DrVeWZomWCOFXm
eaPojfwLfBh3Nf5PDLePniMIGFQZLUNjaVy9xW8h5SPOS7G2/VOfCYWQHwSbt/yw
hASWZUyH3YEJd5txmyYIrHiVi8+GNbr3Tn86BnHRKRbpR27PCIDLPR9v8cXf+9sZ
Ng3JtJu9IGhcX/b4zzDr/7tZ3+DixiO18cfr/Hf07ItS7rgL+czwNSYOmYFduwAL
wxaZS2c7XEwn7j2RPSZIK9DpKlKe/TOD6dYgHbfhbysptQfsrmhIhhqKkhCPoK5C
BAtnklJJnlNMUzk84/CGbJNtmpU2X9dq4uCVou/ZqekqqUhlKSJ1IQoL6lc8k0g1
tG67NjX5O+eVInPnIBH/49chDmOxmf+N6eoPtB3YGQr28K6BDEfrNgt+EAIMGcgJ
/+cptpxT7i3kmLJLIG3yAZ0g+BWgOXJDGSO63r5k6DUobpBMKc05BEA0o5iKlBUo
Yz2/1JFsyT9w+fzdtNtoyzgNsjW/nwGncq6cQLsa5tsSXIeLMgF41oNR/4EJWQ2Y
0EXZ1k8T/7kNuZMs+UEA9oHH/xMXl42qpc2wI7XKHEWpayncHDDE0iCZ2fFCMHbt
2lEIhTIchLKJ4VR8Y4YH5lK2coNYSQp8HS8XK8ZijeXmCBdZyT45f6hfcx3DtMQ5
MQt0HbuRJaXTykAaOeMSw9NjXh9O6e7IbbSOXU81hhJx+Pj0xXg/CDuDvTHMGk4x
AJ6bjCLpdMzz75hhU+WACJtyj8IlFRhqqI4lhSj7KukQcRpLKkb56G49g7kqXyZw
tHSJKCFSYFDFpvndKQ9nIzz89Iq3+/wfY6PNw30ytye3P/S6TtXmZ/5OLRsHOett
Q3Y43hNWFXE/miOWC3bMizqnmf1P3FV21BMdkgb7ApZf42V2DaAMfHEqYMHcezsO
TzaHVQlf7qmjuLXDWYm76xcb7FJctGGKjTBMZUWijdSx1OMxq8lAAiDppvP8TwCK
YMkxmZ/PiY+aUUnrX4zMNQ4WJRfltxSUj56uf3rqDycy2SMNlgA7gs2vMxvT64gT
6an+FJmRmKcGmpZeAoOfFbGQps2mZzXdzCZ8xl8VyoZAzuG0yFH0N6/t31vO3xpu
HtQsi1Bg2TivURZLoIBJPsFyoJT7D8VrBEjyKp6KeCVA1HbLYt31ZlzBaY27cznW
wpxHqUfjJ3qkNVg1MCBXmvSsrSqxLqEyQW1MFONaSzrIXVhrIJQX9nY3qN0gM9Bz
TGh7Hs/voLV3AR+jsoxP/oVIAahTw7DX3aJ0sd//nkljBH8OuStB3PdGXWEdq1gp
FEZkBeZSSOZIRGMd8jf8aFVubPZANcAoeXk5ZWcDssBawCis/4ttDQXgBQaQeCxI
qxSpoi49E/qNeJMM6GdaOZkDSSAy85/MJGwVDnMyjmpPhtKTnapxMNIe6wFkW0nE
k1K8t9k8Skh5eBmDodHSnhU/XYRJfwMx2V2HyCg9sQPg3ZEuNOoEWYJ/B4xbh++J
QkGRp9Y8tUzoGKiZqjfdMOLHVFeZNncVPjG4amgO4pbOs271DyROLWErWGoQGOff
afba4wcpeQ6AQoTfm+cZq/cghOxZlc6LFLNASSygNdDGyfIQMVMnUSZ/l+PRhnIf
2Uo1rC05bzF78DQY7eSQOZzsHB6mGuCTeSePdiuXeW4KMNbcks9Uqqf2gDrbz8iz
gFEElO5kTNFCg7oh3WedBLGf/1RXyY+RG6vCt/Egbf/frjIowgOVVIxLloMSMcmG
jB+USIKy6NAap34Q9tJnHc8fvgfNtHKDO2Ab1p+EdsrPiGwJuxW0anPn62GlS2Ex
pBeC9yneBOyCiF/5P4lAM76qf2Pl5hP+MJlGRYad4lygiSmihcoMBNMGM61dpBru
PeXyBcqcRNhfnhMWsfjVOaOCgXefu7aJpcMFArb4GMYjAbFxcyCfQ2zTtwGAskYn
bUPmHKLpNcz55oiY4MeG1B4oMo1NEguXuac+OMgTiE8Hr60D5bf/7/WfbWEFTqO7
70QMJQp6WxoH6YeWlc9ZKd1qaCo7wDjqAE5sB5wvc3bgPfhTJV9C+NIg1BOqoxwN
C7i9fj08s5rpU5GMRMh8kWViPXNejqCMcZa3RtYSkAKtHj6XsRa1SxzymlVKh+LT
TcsBFIH9OHKzksqQzsZ2nGhlBQjxwQSAemQo82IgYEcJxHFuVpo8rg+bm3+Qj2YD
WtEIOANgqwBYdmTcJuIBW12B/A1xmwgqHbYUDs1yFOQgNTb+CdeW1yukKlPrkpNo
1oBvVFGLgVPeTfHufadrHANOjoLqNrMCjZ557XK6gLoYA8kYrTGJ4Hdux59cjv9i
B6Rogk6GfZc+D6tC2fHZybWiEbZuw4W3AtqFeUFUimNkPjEm2HIYzqX9YUdyTVwm
Zr6TdZxqAE40BpR4GDfRCcq3e0tnwqPkvIRHS4c12a8iu0uBLH4ClNckhaIPF15r
UA4rq951pGw4oA74GVu0dv+oWL7/+70H/9hm/w1Q0Wmn8dsRVyG0DIgfyksOY6kq
7qwUKDxsKN43Xf63FurDB0zn44BBPkzJsL5CdnV9p009zOUbCxUXgQ+eunU6Jq2T
qP74YUjt9xh72NuGQY/KMUYgfRy/GYqxGCQ8rrl2HCMP+/aVfSkhf41KGjIbx0YZ
d75tX6j2yq+8SK1Ra30QufT3joZhZ3D8jdHLbwJvmNilwIFdnXCuNreljgYQ2q2B
FQ70rGslFwORuaunJ1HJjEAcBDcPk6bD0X5Eo/rBL3jp4wVLnOeHfXfX+IZdQ3eN
YY17J+XvkcdF3eV7HF9ygIitRcgk0FG8o/Sdhk30QHohoUU5F8SPYhtwWCYSseBZ
8Z644/YEwYq0LvRL1LeVrRds7W+rFDiDDeQ1+BcE7MJ0nkZ9knyI0/7j86uT7gjf
bO7J2sY+hD1D0b99OnIhCFN9kC5Dsvdo4yWM8NWErPaCOwCkh9H/dxEiRuHHjAT3
GK+L+o2QhnpAJ5gfGTlSK2B4bTgtoprG+UL7aGgIEuvAM/TCYt1w/Yebl7XwfG1D
tY6RtYFEm5VI4NrWtBkujXenMsOTWoyP5EN/C0o5yIRs9hQ+eteSaeCMGqIR/2B3
JGZ4XqFefHbOpyw8D2DNKP7688WRoZcp4REszoJI2FL0l5xTF6eU6fhi7Txq6p1i
T7namhGg3gi2+oA5kUF9C81ic5ioZwBr8Ghw3eJI2me8az/RUboUyCrVSFzSqgjT
k9Jll3yJA4JoKk+t6W8hq/3rubQos/hrTIeP600EbyCO9oxQFh7rwU8PT+LwG5GZ
Z4I/ygDSr2ZLbJeHNg00k8dUdqmhYBWmhjk3IAj20IzRwiEF6fKQpOFS15uySVKh
qC8guDdwAYypgtXMnQeKKR5uep4qOlmm3Drv64+vXXok/D2ucxEMgJWrSsv3MnJp
VgXYIHv2mKMt6F3XRtIEIA2yl0ZK1XiXYeuAE99+YK+KnI5BQJqlcvsUbIaSuTTa
/LjaiX8UVD4DH1fFlKeXoyXvrRTya0i6JLQLyC6H/tJnn0fA9i9rxAPTon4ZEpHK
kYU8zrpPXLlAxjWEme77DsImsNTBhcNMxaiySX0q3M3B5QboCnyQu3ujWrzeCbfK
y/OZ4Uxw9IWHQe1z4/Vc+Wr2GGXjF2joihboEifjI5tXIAlFZBYeOXr0/O/3RFuv
X7JmYei/ntV/dZ4VLKOXdWXH2Od7rxHhe8fMMyxxhk60jZSkl7a+9jq9xvBpKiBQ
J5OJqf0Rm5I2zQtA7sK2/0Nxfxu3oSm9qDSnGvgi+r9l4qL9as9ll/DOl3J32gHG
+fW1AqRSod2YWMQnY/E4R/gmedTVxDkU78ZqzNb8fyR4zEwlwq24246lB7nGQ7QJ
m1+Y/zh17SzgO5CaHjNyFeGCmAGww9SZpkyaA47NJ+LKnakFirVWYBob2F0RMlQC
Bq4D4QwwsWoP+FLz99VGdZ28SHGtIZQiX6acUbHu9oJnYp3eT55UgkOqOUgRG5RI
7qPx4SqkwMtttNl43dtEHJzDxqXiXUB5hw0M95XpmoEpyx5kk63RuvwzJXidunJ3
917v0ns5i9+MQx64pIjD7D7G+BBJ0wRu7bOZEL8wkAEuflBs83WdsVdqs2dFQbgc
RkQZhtE72VlQG75ts37ZsxXHvKVovG/MamiHF/G9c52RXNAcpM7flhZcyOd/SEoa
+AE4w7ltW4rY2w/ERA6MjRgatE3RSqP6vcF6WYhkcusruTOI1sbgkEP6cxgPf9f+
7GHRmsomz3IGDga70lDDEt+t0iGM7wc8dsZJ5rAiASl4H/yDCQKL4IEnDZF9zuYi
Kx/xeHhI+AGO4wIOBJqQDI6GxtKxTbkMvI7EH38dSqoYMo+WX8/k7kP8NfxyBFnN
VHCHlt47oXb3kFO01oLwjGhBy+vZrdABDBLZBx2w0ZoSy/M1gKFTzOqEZuT62rQy
ve+r7pBGvayzbRUC072u9a9Ag2dVETYQ1ZHKWw+mS+gnFowtX1rA0CN5TipeRkZl
g2EOC0G3X7e/Rc417lONm9V8wpTIlmk0ANir+kAKmJbQZ9O2OV8UGm93ofVOLB0E
uMxiEP0UxZMCK1XQYqm548zJQelePQoZ6fkWqiGN6a4mLUl9O+UlQxhw6iLLvdNP
KbHp7CTl12Q781ysXcki/toRGruBMVo3mZIemDIQDXiCFzxUDFik8tk8rVax+moi
cAf2gX0oBSDIFLkentKAmWyY8+L3lt6gsvicvIk+vNGnztoUFpAR8XJYLZF2Zglc
91VKbOxoYLSm3tNIvzUS6Oncq2BX+raLYTieMuoIreV3NvftXIbgaxAI0z9/x5Mn
Yjx3M9fuODw20z+xPPlsnivRuoNkBoUliCEeVDzNAptforBOlA69Tw3bopHVTTTh
Z8D0dIKf/nzh3VgGVqU/WMzF4ONiQNgBW0Dj5N1WjVl59kMwhcOwxh4dJ1qsmTu9
21ZAKMj39x6+/ub5qhYGscssg+fAOgJL6BOEADIgY0/1kKn8LlWnLLriFqSlKdVl
GXbecWQfLF8GcGZbM2iBmSnkb5KB7eZOzoj9Nk7AbXywTnJaiaZH5H9PmOHVt5tB
Hplx5KXb958M+J51uQjfrDUieaZwp9XFBK72gcHhXDbGSfyn4cgGfWy+5Xvjsfqx
GLz2UJIFl1M0WU9In1ZMPXO7b6KKv1+lW1PEzT/1mJaN8ryC8uziQKmQozhilbeN
OmxgILukng//tULOj5fD3UxsKouCQTlFZb4qZL3A+DlQZ47g6cgnndIen1PwVFHo
Hj//ZKLIV8htFTdmWtiET176+C+iNOsJM2dr4mqdcGpIM113AWjTtCQBkE08QZs6
3X8p7VT9fOrYgvFS7PrReiQaSqcJUn4gIovixjgNTcyBT9dqG+1K9oW/DRbUwZm6
iIUYfPci/YOUJaVXzHbBb/QK+9GLVF/SNFoHE6UpfeMcaPnM9ltyzGFE8Zmqvtrj
DGD4Jd6Ikmx2Nd8muI8zRv4YzTDyIf7ig59ZmdaVpON2HRxYnov2nDZiGW1EB4b7
yW4Jid7jIgCWyeXl6eAemhXwSYgZ9PxAG4P70lJK3Hm21vm2raLNdAXCBhio3LLH
u+J8lHSGyP83W9uZdzWPtdFjOyCG861SZYkTJ2MzYGPnsTDiK5unq+52IzmfHL9l
MejMoF8VWLJ52ris69l7FO7WGMmcu15YF9AOqYDLNao35OWMR8vYJMLYd0cCSWJq
83KDKQc89zmS/9EvZStDwWsk8C6ZKKjrxtxz+h3aPTtFYJ80q8AJZvDWP3kpUx9j
joQKa0jL2grx4SPaeNen5HecG2+VvB5YjaM2cACZYVs55y5meBjTYhGQKtUl1b15
v2wpztbQ/udPxN4y8PN2kfrRaR1DgxImzWYckNkOvjEVGpB2B0hF8nEb1bMEFnWa
wNxgdQfyntY70GmiqmzIHS1QVBQoSUglzSU9F94oaSs0sR+FLQcpUNuSYXqW8xZ8
GeLXlUJHU7rSonxDpbhiZsMDHF9CzKR0usmFzr0JL64aSrcPvljK3YOMbkEGOU2s
WsxXlxyUEGygP6DTIXF8ew5ulO5AGTbm9hGWWeFZo6QJ0xWlsAn8LH/72eo/9o4n
5xT5XO0DKOh+XWlX4GiW5amRmEp1OxecJqg4JQAnAYMF3xtWvCBMtQMH4LJa4D4Z
EiMO984CaNbqnKBXfCMv25VGsZkT6yTkN5E92Sbc94mFgECGTVxMayVJXEhz/JmQ
+Q/behsFQnAi56CnQvEWJV0J4XK25uNBS9WTL11o9ocuqdN3XKFjZvkI1RJ8LxDD
qQ2VQlJ1DuXCiAt94Tb9necvINSsX5A6Wc46mOzqOJ82EmclU7cCICrVv8cDFnkf
PhlnOkhlwq/qxs3xTWQrcusdCRU9+wEV4txNb555Rd2IogTfWPQ6WOtOggAp22lE
jMKRsh3M8AfKlqGlvqronuYK3zypgn3BOv4XKSkt39ydaBKIhKTUrfbN21A8q52G
ezIj7Iq5Nww7TMi1q8GyzP2Nst7xA5WoR/mWDC7uVKQyGPVt7SqxymHTPUVvZAAk
5qh3evxQyxWh2SsV1z+3Awg2A3IKp09InXZBmIiM/fUzURIUE22JNVVDMci97jEo
8WIiQCSCtqRIypjUmfRTmZJ0nhnjD2HAPsmVPsqJkEQu0kKm5CTvagzATtLBvVx4
vHYVoHNKrIwU54EljatxaRlMRq3/fs6FcCPcIhgXNftfeNF9PdgtlvrYr3WC+gV1
eLQVncCSgziEPR0sFef3WKYKP1LH9QHulAP8zM5dZMcLroLppSzMAj9KCZ0VUgTY
U8P2GhV/UJJmI5U+tLV99nX9semY1XSajBulypSAvrSEYOaCfbaQfWeSidrr2Puw
SLQRkdhZlKiAV0yo1oiOMZmuM9rY5DoIcftWg1WN9byAjw20vz9Yf+LuON2WiVGk
vbq3ScFIKQwvohmJkQbqinqWwnyPaQK9srCJEfLAQVnmAnVn0sEq3Rc6H1OqyuRl
BIK05gkeOmVR540r7JaKMFaEngwetCNLotMila7tuIQo1p3ZdYfAm3Y+6xXRPN9m
UbBfQuEwpj4pjVePuD7iyhCJ9oWhYIcVyUv6Bwx6pEluzw/hZMjCAwxeDu1MHAoP
mHZXNnC5jOBlyqUo3km2XdP0/47AJXh03287lIau+PJMklPt3WljMA58Qfs8r7jv
g2OXxczeFyPWDdL4EncQAR1V+F5kbj+Ot7UuHrWVACV1NamsGojdMI2y0WbqSUsW
qEBseU7Cjyr1MKfQqKE7NE0jmVPS7ELCRfBi0JPA5AkTMO3han/YWAihQS/9c8eJ
FVc3fQ8I2OQUBEeQ4x46tY//v254fqI5/lzcs/7O5SvRoIatRoH34wr4EH5+U2Ls
cs6hGWHZPn0Ajv34I2wvP/6t4rdRrqLaDUi1nmb5B6LQ5eDxAe+qEw6Gb0d2xMrv
jg7QvkKRnGUCT21QCxGYxyzqq//KM2MrcEd/HjU0QaClEg7RJU4l6ARZJavwWUWX
9lAx3ZiKHUHENyeDMCQmEn4zSVXr7pNKoARqeVPvahGInaRfmwx7WZXYnWopU2Id
bIX8rKdU8IdDkeyofH19a7KFrJzslD7brVjDLd5djkGlzhQWXxT/BSyXRg8kYLoK
/h35CmPMjoDMZfhIMbJw7EVLO8TjIH4H2Mirf37x253KcHfvEy13+w3xq5wn6IV4
hgztbUorRUcBQnx84VmhVLhf3Hygb4giaTtDDZSQM/DxhpFh1KdOMaGezxV2mEW0
LZ7MmbQspoYHtABLQMgvjTmp13UuBi/iX/FJFQCKjdlQkePF4Aux3GBnMDttVwZL
HKx1PC53MxFs575RabO/DBUmo6cZwYozRiSb/i/O6h+GRY9UaFOngqC7ZRoXDvjb
xvBUOANqRvP9/596xGTTil8LYfJtMcgDBf94gnCEkEsG3KA3ZG13NqOUS6eGB6GS
j8P/9oZcoCFJapjL3I+DCxS5sAMMmfvGpq2TJ372CQvQEj6Qkl7BvykzyU/0jEw4
pTBVjW+gHyk+sjV3UA05NXvxktQE8mKgoCIspLkQQ3LmRc1ktEB9LFy4w8HAPJk4
kj/6N1VvTVCNcJwwqYFKr28FIERuKeSTcsOahWoUGqJHwr2YjQQNhpEAkH7GMMzF
d/qRRFYJPNZpKeZu8YdIYLn90y+7kApLMwsrEtDQxYp5hZe7LY0541lw552Hf26N
84IARM43SeiXXHootfyDtIZtp1p0haTn1kfc0ikZCH1KKktBMXtcjhHh50iFjREh
i2JVYI611vxDeCJEVI7VhRQvXny+bbYmsGXCzjXNEQCjeqpqoorQdgJbqYq3lhll
+dp/1H2/J2u53MGFCkt2zkUubA45HYgcvW6lasdEQTcKgLwI+sM4pfGZI+0E1ZJt
4HCjAoFY4QWuNyFWXsPnRCGDFe3DOuiJekaLIvUcLcJXxxG0fQAzyXdfb4d3JeNo
rwuArVCy4pgEV7eR/E7BhX7PKgKRMUMc/Q4YjAoxyaOjbS4P2BEK0nHwf3LSEKQL
cSq93Pzxdc0NPdnH5e0sXwOz3uy2Pq4xANT2Q3CL3WO8fMwF+b1JNMMNjtGTl0Yz
Yh0XBTt4B8/Av6axmKDJKim2FXIZ66psFi0wbEftljP+TvsJTcFUeTknXIkfIY/u
ridq4nig96IkMv19VXQt2KsAk7K3vx48cfww7bRyYXUeKyT/TPf4Xjdyx1ypV5O8
PPfP7mzxygnTjI/G4ZoJrzOMv1FrsPB7NchZ0bfEorYnyhlJIqtLBlnnm9eiza6P
jhVO6L+4R4Yvz8MKyOHQPZEERmyUe5gp5QoCQ2bRblAisRPGtEqwTkgnQ9BgheNj
FnrFjcq1xAGEnOW8+qKrVjpWh7iUVf2GSvkJw5amUh11qenkERq8dR0uSjNAf7a9
QHEoLmuTSOFYXurblv4t6tYPgIZJ2r9akfsahTOEaHaZDNLV8SYt6iWGOqNrhYGf
kWjy2AzXXuXTvVJYm/QGmXdXLwhpezxB/cV6fFgHonAgEhWeQM9vZszuIb+apZY8
KT2XTAt23NrsHRymqGYp/VRt0wGy0LvW60F6t1fiHqFyuxcmNkuIdb/X6ft7pByL
o73gqIN1sgmPPaoDyJN/ZLYnhZV1w+bbX2NMvtDq7YHwMgDdsZ4hVkH+jGHK9Vc+
tPHDkcxeEapPc00U3w0esYlyodgBDA5j6nBYctC5h0Ryxqc3/LGFIe7lRG8xzfVt
vU7SjjorjsWiswoKhx9hcMoJGj9w9fvCNca+UO5I5y2ZaVsirrD5P3XsPovzTQKn
ddRFP/HBf1AA6yjb7zUwFAf/meSyjT4aAp9wB0tz9BJ1TZMsV52S8jy3EmCzWQqS
n/H7UsZ0wGsbmPzD/WF/9NmU5/9Eps9KYSoWDvRc/LKuvy9QgN2jJMwwuW86mhSl
n3UuSBHJoJK59f96wVXkuDOLYhXIxM28p0NXUeda+oDp+P88RWxXgFYo4cSepsDm
i2CPH3F2+uNv1755jhPXcbEdDRF9yu3dBuOg+4l6/6TZgolIWbMjAjYv0rAurG4M
cRONuLJN4h/mUwVsmtoAP5FKHDD6pG0rJt7dIo8h7n77Y2Yui3z5bNUF+6TID/gt
5Wj84Pp7s5HgFg7/chx7pN/ejUWC1R4slyyyrVoCUubHYzYHlUtrR+Ldy1VUKnvn
zCnDr9J8U8QGx0C5b8u/eleA7aUSH74yHXFvsv6dJ2vJpZ2d2Yw9Leh4swhIExxx
G6QX66ECGfu9GrogljJXuJdzPR20OAIljJZUBgEiP8+wlxa58an2uf1gxxzFeiSZ
QN6wO/1jinB6AZLYP5paSi3Tb11I4q+8Ah3kUonYp13AIVUHvBQF9FzngA386qmq
4EfqYxYFKrmg4YIJWRT6LOKcr5zFm6/5oVbZL0lJq8X8MW1Y1tatdp+ZPmBgxb3v
T5HKD1Rb2zRRpItO0YL678JhGFWoREoFn4FGuUUybYs+piYoUqKfsVdxHXWfrlDh
5fHTGzKSiyVjj+VDHzp9VhI1c+r2G6y8RGw8Kn7P/fw17/hVJZml40j2RUNEQcx6
k5QVfi2KzJRmYZaCj+TvjVZjNNlGSNEuKI9lZnaaFfzvThTm785t/q40DXdhylr9
4Vi+JFI0MXS/oqgOKVE4ozZ+qMvVz25U1jUYp6BoazIllPd37LyebbjJT9ybqGs1
UKlN5pHiOAa0Ux+4qgEN4LQ3pHoNQ9tav+jgU3Tuf4mAeKdqKk71zPgwEDc+0T+h
0ff3zoN66+XbZG23KrXJ5FcVlao6J6RqBYF0j6UmdwDa4LRJB1DTZ4PPfyj5rIAk
sfR+pXnbiDb3044MZfYHh8Af0rAM1zk105fOcaNQBdKnGFFyWvjyfqmUxj8CqaH2
yjxk9X6giqUp9GbtFCXEmwIa9OXvHHolSpS20956edo41NNxWRMTEAjJjq9EfjW5
14sOq4xEPhPrSTzDrE31xHsUscCedmuImpuajq7GdvZxW83zWDStYUrsOik6WukC
PYSvBehmo3AnrOyCbhNxownz5YI1aZkNfNYPLP8IqKRvb+/AaAbHmSQDUb1Mg6/m
Po1mzwI8awEiQ4Boq+KyFbYcvk1Tu+GGYkKdS6YHSDWSDBBjSjNmjr1AV7pOiCHH
kknlbkdLVW97xbwObJ0KkpTWpARQZPR4drBNM5GEl+16NkxtHcgNWirzC3F8vtEl
UVIbLQPBZxWsvuMwH6CjW2YouGlS0ovt8pDJCq9fsSqu9IfkSInOEdzo3gqhmcjt
Flm3b7k3EPNd4ehf96QwLFdLTwHwzikS35YY1rDXD3L86hQJ8brKEeiPCpjPVV8y
UI5eWI+h7hR/jbFGEM8diEryDtBlHOzdJi6LHMdMDP6cLP5Y/1OxVShF5//ghFLg
Tq79WfdddabxWdiWp7nmOvFnttSs3kszOdGLp1l9f+PHAPtO1jiSPR8BF1s1X7aQ
CaYNDxYAYblj/+ECbnzAjsTesMtcVkbLm6pCk4lBMOIqkW5+sPb/pg87n9tKLmmm
IWC/wAh2pu5d7r07RdJsAAyuyS28d6abghbOmc3L1qAOdhcBO0jeOS9TxSJKLmHJ
SDt23z1ivzQEsGpWjj3xw7e4nYj5p89/puTgUjakANmOnK4gd4xiXhCtxn/nEbhb
D/fLzg3ywGgcSU4KesAnA1DXbrIkXGBDVF+OvrzKV+uK+nLH1r4zFv42ZFdz/QwZ
cBWfZcpaq6t+Pcn6iYEKvn487oy1uEhk5fK8cmF/DuzcSm2jltbx8ubQb127Hdex
G5i80+VIG9MxuD2f+BqBKPoDoOFEeWwbQ4p2RKdkN6nj2PIWVletuvSRgVGlwD3M
kOusMVAt120njv0xy3HxNprxcSapxtsh01D40LcFj6b4hfzqfuMvPZlUhcOj49eK
KzLaFJzKdvcGTYleCjxG4vizkiqcznTPl3jTyPDxWCLQ86df4MbFDG5Zzv/XNTWn
od65P72j7CCUjmzKpupanf2Qvid2xEu7rzF9+JmZ1lqOLL37BaLe9NzefAuSBD2B
y1mDPntI7jPAbxBRcXp+8h9K7oTRgI+9hyqg6TupiNpzs4flz1rhQX+YSOaJhSeC
QvEQSkpuqHZqKDz3cD5Mcbn9tD3gvmGvtvu99vbFpwkB+BT2XTN3xyRSwAbn6zle
R+av7G/j/wYbfc8MRonpyxtYUrO/FMK1iIpJcFRTzHRtrbCyRq6XGMjD3D62z3SH
WO3/QQLRvarTr6oYaisZu2ckIBr6KtMgJpb+WpybSXrTcZnwCy/PGB1JrIl6heV5
evyJSYNaQ1SKPQXpwLmzLKM2gLxpF8gXju3qqnuT8niY2zOc4b7c+qsj8Vwjnbr0
+GHqCo2tPiqPnCwU0lxN5d8liWdxad4iaVzDkuBj83lvp208CoKZ3bCWBh5qJoD/
LXvYc3C8xEFCU77BLx3QHzMDiSxsdPIeIPU9kPajXjxS4qjVyMbDrkFmV89N2Jtc
bGKAwR30crX25lcJDqTBVs3U/Iz7OObolqGdTFNexY93OEvoTCJfC2aMGO1tgLJi
13ZXP8a4xq5v5rlTZWUO7XJawv8c1DLnyKXiOMKUVYMdEPcQ309WeRvaT77moqgB
fCUM94nB2ffL/vMgKASPBanPZBapS4sbpZf6LpimrTXDMIIo8ijrjv5DxOO37Ly5
NXBOb9U2VnChd7iUF9Uzkd0KKJIwaK426WwsNEsZ3wbfDKjMA1prN1+TIMiGuiVf
6h8kN/5kcTLl2lR4c8KN3P5QcCvKLz1f0Yy65YM7MTO3qXJr8XIBf1hSRd/CDAUP
KmAFfMbpisweJBt7BhsVlCf57Kx8VeBEbV+wcs6CYfTvsGJAw6gEJqHmAHcaQayt
ac7BkJXSuJjZ8OK8CthdcHXlEQjFNEc7s5sbLAsvxnfI3KLje3GVhfhbEyaPU9my
kEFnjabJVk31fVqkDOMV9dwR9ijj3NrrRF/zV5sNwqdfDq1EjWe/WXkheWAWWQES
Pd9Mlv4eB6JiZklcjrxn+XF3Ilss0AqIux7TPfA4i92emJhkmCQTefE3/cp6PLbR
oZe7+v1XMJhX6Jt67o4UmmhxVCrz45vmisikriP+CjHB8JuZoqirpqMwWg2QWQjn
b13e96N0madpdyrxe5CXXufV78ocK7wGSFlPD9j3CHpKwyou4H/qihGXw+YnW7dj
Uh6viAENbkjV2DmMcQVy4nZ45RrUu92ZpQF+nnlxT9KKp/no/pNaz/07BYIr5R8w
1Tb6MI71iGVthluWYXgslulNx1kU1hsrBzt7gO5pGvnOONI4zYssPoKDpsYhDPu7
ngxTj3mgrcWLMcYE7rLfQ7Dh16eUXCLeliGIETNW5zgmXY0GlImryAAdA9K7SiOJ
qMXHH6E08rCetGFxFNQR5G5ErJr0Hnstqrhm4H+BQtiCwAaJTJuOVikkNAA5gBJo
0MyWjPXFvQXN1w7aLjJNPGkkM0Jc4I20R9SxdpMV2BIm8rCtoCYTE1u5+TpIesYa
v/8EqBkH/a/lKmmLCYpbK6rGWKwVzSMu9UyNs3fQJdavFXkHPT4xyDcHHhmwN4sh
vCYQmelT8LwWnJOXGsdoPZx61SD0KbfG1ajF3ouRc+GjBfoM7s1l02lDILsy501J
GRZlbZuzMSqNX27P613nfp6TY30OHz4yfzCjm3ORgaDeDXXwRBYT/OifuQ1UL8fK
+g09R6fCBSSbR9oldyD43HbbLZhxvN//p3/Ady1Ce5U9Jrt5N4XnT1Lcy+hLPCfd
Qm219VxC0o7j4n5ymM4W0DfmIR/p7J6hpdUreo5i4KcMzOqTBZ4+oMOuovG77SsW
TGtTvx0M3bMGmvxfwFok3VMk5jnqk4iRRbwM+j64BeFWu0V7Y8vl25njOKiv+xmS
2IQute52WhACwACVib31jNTH04DPu9Oc+SrcasixBcyK4kkOVGaNVMuHDDU3kBPH
kz3PC0h2Ag7Gmj2n9AoKuduQ5JLAMx2Bubn37zEfMaQ2OE7tvOQzyVzqmRp8XsKx
16DpoxIwUw2EsQFyK6ZvvuMkNCoD4UjyvpiStJs0YP8gv++XO2e6fAPN0XQRRga0
le7P1NcsT9gfqYcEDYPlEoGtnFoBdXyYuP/CRsZ1H3YNMqadokYgMxgH3+kcGC26
bQ5wVguJDKEhP/GuGNQGlI64IOxUsFqoHIJOetAGyLl+iFH6g/hv0wZTffnwR9V9
9PsfX6v11jK7tKCXWQ45f36YcJjEg0PtFpl6h7bjZ8X0LG68rb8KP7g1rAuIPTDN
Bmz2H+0zAy90eAswVOksKkmoRAq1w3IC/M8AzrjJhl1wygunWQC7vjkung8FolLN
epjxg0jI/9cC0qlv4m3LCxvfYw6K1mZubZsrpboB7OwnpMCXEFkUd/loIG3L1CF4
LUOqjIGmgxceYl5l9KSFfvq3m3DJjz1X88sU5trrT7A4lzwNU2CAiiQV4JGjTh0K
sum6JbLOi9f+JXFE8zqoZxkIrxLaSgoMYTKTRQSsR+bT1f7sJb5R/D7sDOJCYCpS
NgQXnpEVXUzy/Kekpc/5pwDvb2/VyL/dN0CqhhqDr9Y0UXjlS1lDZcwXNUr6W9Cg
9GE0JSWsjHtL1Ti8R5OgxjgLbnZM+GFOoQ/+Qpv5HPWe6H+mCSyRo7ZI7d2ez09p
gBuVLx+AC8F2M8halSIzJWSKQ0G5U/AyBC9oxc8HnludFaeklYiIyMEZP8pky/Ns
TmMfyj89pTQkogykk5Kdfynu7oZp0wGWis+8UWMF/xZfxVfrtLA1jf1nx3OeQjim
D5N2vKD0Tnm4qH4rxMxwNaHrCn6oxmLrd5WQCpLDzmZQxTqrDNUPla9+YdFWgCen
y1iRIba/f/3B7R88Z2FlyUCm2hSgSditrEe8wQ38dYbfki0dXQLXX65UmPZ0Ut9J
Bu+3RJPPd/lt63zZIsGVJtZmH/qhc2m0jucXf5aU7f745SXcRJiNKSCkgisvSWpP
ZTHnAoYcHYFVfdwRK4UK3DNfD3msH7yknkF45YiLQQh9b62CXAHyMIrLoWIKwGsH
km4sOHrgJOyf+gMR6OY04MbjYFMPZTki3ODjAWVhYFLteNGxDLmNd5dgsxj6LdWk
1CqEwa/f0W7C3SntNKRVdV8OuP1wL4LttC17LRPRhNrJ5ToRLLoDgsoWA+/hy6vU
PcgvQeCZv6lSp6JBi5TuZdZ8OQWTp3c/L4cCKjhXELfREXRiqfLuew25HSAD9y10
BN1DirNpTTkNIP2gdzAkig==
`pragma protect end_protected
