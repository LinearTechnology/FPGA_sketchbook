// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SWHzLA9UWAKPfG3YNd4oRHM+pbd9sovRLV6tJ9u9RxaRbfmrLvhPCNgTGAqVAtgF
/C374O9VsWTP/sZXIxRIg7sitnEBqSpvL9Hikrdk0PU2XJJ/T/ASv2yofUwu1bOX
4/6OAHWHkWSQvwg4ioBmGXfeIUPxkBmUaTDK2hFZVmU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5632)
Fg1YEQDmj83dHfQGO9C1NQarG0u2PtzclaoVLNhAmzjgu8RdoWgwxuEqiOYB5sn4
FahR/qTQFe2DGI5LQrgAepXwSiia8omU32/MS9FyePPpdWkuzeA3hjVSE7CTZEdR
FqdFqoaMI97plPOXf0vP8eI832K3iHVLSM8gzyOjvfW1h9ipI3CiYzqCUVLopEq5
o8/O6eYyRr6VjRJQtD0OTVOyCTzl+kGBuKRSecdH432SzYrugXAXofYPAmcZ36NS
lM5nF6PvxTJ9kzcvmGgD2xpIbGTN1zfmiGeqmMsNRgWujPVmoF9gQPADTnQDaumS
Qd2PtwxlObJHhCv4jb4fXiw3V2Ia1FSd64/4WEmefyhRRZpVVr4AMKL9cvBtl6I+
vPx2dST8jvgN0n6h5FRwB+d75YOt8iM1n0kRc6F1OPCk3NxRvWfyizrua+WdExl1
n1Wb+VXBQAgsixSoeDQwVNdc/C86nTfXMOx6MMK3S8cuhPRkbeTqnlLHvIq90IrR
/OunIWEv7T6ovPtDu7K3W/qP7evpdBcZC5bJ4xBSF9Id39OYGJbdtcI52vyHBMJF
+v/klq64bUN1hphfbpuU/Pc1YOkHJbQo/rsCAdkUFYvXbUPfxoWPPXvQodLrpsm+
zXNa4Nc4awwf6pBy6wWb2JE9K3T4I+4yOxiB0U09alfpWTgQPeUpxed97a+tvCVu
M059CTyk8H54qvVvPvTXHvcu/zEIUYfHBKgGbVYo2P8l7YebaoqEUgzpqAwkwqX2
32eHzstBQSCPiAN22Wbp/GBZ0yNw1x+4KjvjRdXgZjggF9SNO3lzu5p8WqlIZVUA
JZa51wq8XJPfuT9u59QWNQKaiNm7rSvixZ0EKvYljwW8dlkp16W1q+9XwnRiMlQ5
uNKQup7j4NFLW8MnbQr9C+t0lIkiu3PuCZ1XvHxXGNREpxbwNVAvfH7Gb3MtoF6A
VP8a8sNrcpEoEj7mJ4cTkvX/6gsVTGE2Zq1XOd9kpu0O4cqxerr7jrxsMWJJouuE
8C2pljPYatOccp3LWGrY/KXo2ovb7uatG5ozaPIoECOT4X7uTAZSUCi8xlbedwdq
3l+4NLWJFVU9+KS91c3V3iC4wM9ukLnhiD1JYAU/hjgFZZ7pNZNZUAp2+KsNOZVL
Mp7YKbUIlCDFo6s/1y2Nnl/5OAXXrHJ9o2bCW1ifDQ7QEw3GfenAf9hvlQO4/68R
6opgO8GoTf8Z5tHU316mdaBNzIYKNmZjl+ZqLinFWhKqlTQxKhp2iLGNKOpHsD7X
/OvgKeU9RYc3/Co8qtOdRMo1+YLafQAz+wLxqXex6/p6pH1CGo7tZ/GARD4azZgF
VlN6dq4z8h/0Dg3rLVtWXHQqhIXl7GI83IVZaYiulukC9ZJmiIg4hi0uyouvKjDl
lvk35TqavRC/TVd/8UNAGQ8w31ULCKeXSuB6ykHl2ytA7AUB46C8DJPUMOlF51RB
iUpLZf20V0zm88SMPDSrRF2AnGyrjyx09DdsIJ4raSho17ZhCOVE24RKpwA95DHh
mG3SK2O4fuOgbMWMmFueLzwEf6GL01YvusCFyivauzaqdT2qOz/Ed1O/ZBm6Jpff
Ziqgv+d+gg9KkRxciFwbzUkONi84J8Pgtq8Jeeafj1mcVpYHa+4Ctaw33XNuNsUC
1nkQ+a/NeTQknukbYCAxTSfdRbtgqpy/W9wPSeuApdpuAk+g0LlOJIi+DT9svQ4T
aW1gjU2avUX8MgHSpXnR329AnLMNFq0i9tBtZJZOq4DQhMSHeB2SjGWENTlMz3sZ
I6/c5biGmfeUtCtdhAwXF18kHZV6M00gIiTKSxvOke8EE8Dt6d5rDKSlavfHt24b
P3CYWi9H65X8Mr2cweT2SztxNVDMdyvmjKhnM9HKD41VWrr9jnfRPZI4vCaQF0CP
E4VYI8A/SNS3kDVrD206fJNwvdKxfxexKjUf50uA8USILBPrbgqY4SJz0DPhjfb/
DcTW5CJ/1DocOhcnJR+7FJT9yvCCUesvlUe85k1Gss3cCTPDXtUz1wogaCTby9ke
h6W3C+m7bz03V5oRKOcjsRUcv3I929pkihdEtyMFdzgp+F6YNGhVY8tYg+vWQ7Ke
3KklAaIJtZtFc1VNIo9OB/hoRbQvK2deJEIAuadNPnPBc5VguWZ2vAHuiA8VfE5g
rI81FwFZ7pSWdWAM0i2a313h5VlS6UWylyWKYxJdjLicLAhdGar1dKzkRfU5LX/5
Sr6MFa61Hk4DmSbJg1SEHsMn8lfr9pjJ4NBV/hdpyXVTS+EFycVwWokw57vGMAia
HDfY147qhTLsvCvjv6wJy7h2OOw4oFn24uny/F2sYvx8rvy36DZS92ABym2q1KmZ
//PVH1RxVQtoMTJ/3owKF5ICwTP+/kITolSnUUUdtTuvMJavmFCHQsT5dph+7R0C
wj+vGdnns9I7VSChwaI+Jol1y4eD/az55D52R+EInTpsVWPW1GA1GJpRL0uaB1yo
mB4jR6wN5HweYEJgkTtXoBTb6N74FREI6QW6P/xTF30ErwfemUX3I8vd+Pe71yXW
fe01hROGMjlQUABrC3Fqsx1HTSWHk0FPKaS9nrasb7P/xFTpp2MNLHZVDhdqOqEh
nY8YZgrIfMK4a6JlcJWTplh9Ij8yolIzh9LFGMAeyy8b0c+eHbw/wrqC+2+WzyFd
TKn4I6i7MrzOWuR3iH9XJ1ArkWu40J3SToggnA1H2+GnylmB2ACj5ZbrsSzDZlre
Xn5GY71Qvn8ZfCil5VyTXd54JCxjF5zp2feGe0Y8xfo6lmwQkwwJOMLA6al/tRRR
BhZIVPb74NKJ40j3qUnP1Y0bpl1xrPuRS9Y3pfhplHQe9Let1+cWFJNRWi18/tXN
ldExWHYgziauNUY6M+EPcm65SiBoLBUpjicYXJ4oxPMqUNfQhnExP7BEuWiuc48R
xqVhvTH3SbnX/Ol1UZK86z7MMJ2YqGIRwi9i46S4367zffemacK0xvspQzraQbA4
3QI8+9x1q2SLDVE7vDJ3DkA/S0ON9HhcB7FaSWHS1eIGDhEbeIiXTcUUr+vXA+ou
HxN99ikBe6nLPx65NrZY8am+Fgpo3/kk7ODTc/Z69kuJN0ho+QNlDFUWamaf6Nry
7RdC0EFv2S+po2ahkdpEkMlAlcL/MWYFN+CnXJy2olHZ7A3iiXZEr+b4X0oZTwGk
By41j/a74W1UG1jUmXIDf8xu+hWuEX83wXojXEPj/gT3ujQg/heTtsyNXB2ihFgi
EP6Mm8f09cIy3KbY9RNM1auHwPrQniPhXrOnjvkqqk0WuTesGJi2xNTkuOHOh+Ij
I820fAmjs6UrQ5m2SGAUBpm/FszEz7gkk7WL8/WeyY7fKObAx1twQMyBzFj8b/Zg
8FA5EYBJpjD2n3CNBPZbbgmxdWzfMNLT2uxj9QGFHORcgC0DruDiVRUei2h3PoWw
4hmMxwKwx4RvvPZtw8ANDG0NBX6mSsJsMweSbzxqLSCLsBoD/MfsAdnfoKLwg37h
aQNW2cZmgIOvIvY1lw+Wv5E0joBHBh9bc2E6NUsXigoP+qZjVYUhHSN3YuL0K0wD
GvcdVa9A8BewZI1lwkb6BcM+x3JYb9Zd14/m+iGwQCYvpUh4vFA+qNb/zUY+ZvRV
Y5fuhYfRVKnEZMP2cF2R8RIrsp6uGwiDEnA+4a02394WGYV/zYArsfwshzgBVRrQ
ymIqxRMfXStuqWT6pLGQ58HCHhKGQUhBxEcKb9rR6DXjVubrXgqtDTEtU378s5vY
jJfnDMhX802VesgVR3lrKSjA6SV/XxlBX2QrF7JuRtU8bXglsCfFsjeDQBiHtBn7
i3G9bfrG7HNPxGahUFVwkhIGyH3/Ah2eC9w+JN+klVt/pplfr9JcK244UtBYn/0M
uzi+uBCKgezIGw7ZtfM3Bu6ZtZ11f63Rqh481VWX+0xBocRok2JmlUcWgrCV1vT/
lZlmrEQRGd/vxsPh+AYG+CM4845j8QyO1w4SYN1kK8uWGrLY7dHyc6oHP7gEGXoQ
qk/4gn6BA6X+K4iI4AJrMqTJd1qPBLk2KB3oIjJBt5PIPx78pY86FGV8F9oWo80A
Bg9ZcSj2R1E6ZH/llYIHO/pak4fAXOEZjBp02IgOFp3jT28100uMkIgc4drpJ1H8
tXraJGlkUZSO3ME+JizkIYvMXdrRqL73X6g9mcyuOo+UKac9QgAR7gZlZoArbs+v
lTpfBQZ2Ltdf3jbcfVEeFnvGsNsKmVbjkdpoULDoZy8XF3e84w1J7wFVCXoS13vq
7FAYAkDHhKQG/rYxaAZR+BIgRL0ccfjNLXDg27HhvLwCqSjuufmig77jWHRGkA08
8/lNkqzH6R1E6jNgFTqlbLwP+bmfigYSL/Cz+YlerytQRNx+t98zhGuvWlPbvv5y
RYMhc9tmHDgJVCTKHVZuBg7rzUBPZHXrCIj0HK7P/x6+wEcwRs47WT3Wp9mcBHRN
9FNd00B+iXtQkfWW3nEoGe2PgST0UxMJ+W922+YOwvMKDH4ak0qwvhAQWARi2YG6
nuUI5FbZMnVF4LAI79oFw9Q63+rl+atnCm4copFZHFJAQBZXMsljkOpRLxEUsxPq
Bdbb+NadBvlln/Fd99r8XW/JVSzfp6RLdXcaWTrAuvzVfoiOIVSkBx4+dRymlFww
lnsxoxuOtoO9/IUh9jqZhc2suGkBztSjNGu70EaqyRSIUljOY6gyJ4u7ajoQobPC
YK+aMNEzDUrXYwrjmBGs9f1oHc/9pxka4Ru1fkTLkgL8TXwzmmlht3U9E0RpBnNF
O+lrb39AoOqx3VldI/3nWGqtCwvXkL6ZZCTDJk5bVio7oSfFRSVlRXa9GF/PcP4C
2joqNuWnuBN8nLjVhcJPLCwHNRXRmT3ZZHjasI5k2UktWu06qZ5DvY4BpnlfDIvy
NabvGPSYHVtSlt0+m6ar5iEKW535R1U7aGSFtkEwNHxH7Gzeo/7OMTX671FNdSik
Lz/1QQKfapoFyz/2z2jMpOU6uhbO2AP/aSuC+ycraCakMufQ2gt/1w0sQgFg2mr9
SSHEdHHMFeeLfyHwF4PIVTU/PMKEzBZ9VjyKpCx/KRWAsWbpVuyjMp6YxTGGYpeA
OBjMcfgw4pDOm1wy/ofMq0tVNWJTm/IWE4Tm+x0qVYKhiNOP0P9jluS9xdjVf5Vp
I/9Hz1mGJVY3kdSuXHpCD59AFZZkIwMiSDlbiE6zCnNFRy5vVNEmNCvjQ+vAedeU
etmKB7kGClFn25exAa6EE6VhLBMrv/5RPVSjX/JE2AyuHyoDSd6cc80utxixvvHk
amK3BlZAUR1sqX3E6v4J4eqRwLMsAabjlVJo7MLkUE+z6dxc63IA49fl4dlFnaGc
Z5EFrZglbP/55jVRALHGB/1F5uhdewJ7aT4BS5LATkPH6uqpYZSi6JxOUqrHNdzy
ZRch7Wk2IEBkOlghjh24BMxupd79JbXTYxeYEEZWTIHsXTCh2M+RYFEdWiBoFEwO
qwAoQWI1p0SPJ3tkw8FotrX9wtqggXJQmKLsVCQHV+Yo3TO9GxXzyLBHcMdSA5nq
eDashMpmUJOpWH2yWDgiQx+eb6upw/Tz16ZYIakjNHx5+qYlj+a9eNnGgIfuClza
r2c0JATLRSU6zG0DWDaE6Zuby42cCwDD0Evl1MTXh/jQHc7PGp35UDWUSzt1Hgx8
19vmi6ulnJsEWnV+vv27kiunutklxT/RFqVAEiD4nEZ0Y54Nao6Xj6Gtv+yVruzF
9VCVvVidm+77NCWodQjJnZUVHI8pJ6LjmE8LeJfIpgyomKMGnHuyswT/240ZWdTW
3kSRbZnLQyNjrXmpZmMWr1WGgvQFaQRrA1fbcZZ9aLSkK6MzAfXiTNRMzdy3XTLp
eaxj7JBioscxQpIFk9LRRXVvA4BcSki8/FbMAWU5dJ3Ae54uiGbtXuyggOTJuL6d
S0iNK+YMFLVYypd58FioE4GCTCIU9QOqzWOKxcKl8NZdLwvHr+BYasG6rx7ECQZH
fFN8/cKjRxvzL9FZ8neu0h2wKEqYSVk1w6qTpmqidtYXNIu49z2EHIDb4lNSCCok
bxZjd3joYt2dr0MErztAanKQGenkXe1w98pHNikDxduM3cpYew6DmtnOBZTVy+qp
M7U7SqcjmhhkcCRf5zDkLpA02yTse869Oc4H/7Lh5VMDamamhCt/z/d48k92KoPG
jFGSOy1AuVA+ImxmE1gkgM+NkTYtg9tRAkQYj0ogU8yXwAuwoy7nP4rFDV5I10xo
3WM5AorlZc6MUy06Ly62lPHc2rADZhAsP8+I8zMlAP9qcp8u2bls+W6dFKhHbqDP
1npLckrP4S8MFi2xwA0F/80PxdH2QlIDXlj7c9rzvtJ2dooVEr+oxyv7XYHDfTt4
HqjFP5beohimPj9jMDBOiPP88ovpXz3SEdvqRTOe4UmMvABOHR1l5aXr1rxIY2V2
y4PwRc1ywxOiPgX6JcMmlhqH6n8Jl6qj2WMA1JRuZQBgAm4gWn4iM1HAEer1oeDi
azbyBO9RSj1Y61NgytHgBPTQRIHorIO2Li/qfKm2dZ1N1cDV73TZiribusZ4bovg
uBv+Mqf+lZKWA3hKb/N96l+vk0D2xzdtLTrEb36atujRbOW9j5G5z/hJ0W55AiNz
NbZZIfoT7asak6Te8t7T8dIwJojOhZEH4+p5jUb5f5Ck++jCS/PQSmB3tX0w1w5t
AcDoShe10LYc0ydHNy4PTX+JdRvVafypH83bzu0TKRfoY42qEPXjKKDKj7RVGGsT
fwUzid/naNYk00dNG5HOIMJYiIYt5qg/neAOI4TVbL7M27tj3yV4dM3NG7uryE9a
g95A86HK0OaUPwPwCpmi0H7QfzSO3otFpGGzHPvqQOZBivTwfUbW/k3VaiifO3Ze
xEFp/oXyJPF0H4x+xRXYk2GGwRuLm8ZCPLBAgGDxlsY6PrXUi8SDw/jcSU8+DzOk
tDC4sUCeLweREstdPrtk7CyPyYrteGOBrN2UW+eC/jcFLEeqYqOPmmtKw+QQJZRO
vhhRpoWUqn+uaQb7+2a/y4HAt/kSYy4KE55+vcxy6whBY+lFsThtRkfvQ0tOVwmT
MQmUyK2++8Ocz6wUAEVIQmxqhU4ktCgmqpwDcN1djQs1QoXcnbw2E8BYjej9qvZI
MHyi5LhsZLEDc/s9GINkoUvs6Y3AfmrltSlZ4qbdboD+zgyc9BnoqOXuw/oAdEnv
ga+5MMxLuZ0/UIJOfdrk56TJl2qhyiIfSEArqo+b/q9DIK9r43WYobaHepOz2a1p
pZ1ySkM2BO1GPgffWaQyTEiMlnGJ7tVsZ3zYUoYdhd8Uq0IbAkm5yd95QVjMndlK
rigR02vaC/hGuAWnFY88Cwu44rJg/qA1lDClA9/186NHb9OchHgmhPL/2eErTwQL
rQ5mfe7QsR+qCE0NSLz4XEKZnBLiqoGBu9Na+vD8+KDAhdnr/vMIbefOXYyEn9Us
lfZkMKmWHw/LSlOcP+f75g==
`pragma protect end_protected
