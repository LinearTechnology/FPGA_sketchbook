// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:08:00 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QhIG/CNCSCC5Lcr/rnLTtoEbgjNkB74NVoaQOyY7DQDiH/Yhf8ZZmJruow2f4ukH
ZepXlrgZtZh4zBaCvUfApPy9J1YI2fXAMm7QPrbngyCY4TpIFtwm3s/QI9A0Upxq
pSXOqXIvolgWithwHnuUmKBwkGKXH76TDwAwAz+2Eoc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15744)
1tyOP1Xrx2tJDQkKPbmqfS9Wie4j+H39BatWpaDfvCQrFPO3leb76fdeyfJun++9
seKvj2D64+/o0GNfZ3QktEGlWP/DTKuq4n3G9m12q8s+ZjHTpt9Zx55P6X2yHRuH
wz5ngwl3BUfA6XkLNTxa+5dC8oLepVrm94QiD36G/sW/Jg8PakMWsN3YkUP7DKth
MIqvl90OmEvDhUGjgc1yw0Gl4ShhvqXOXOI2yYzPciBvYX/eI0K7IZ7uCWu0dxUj
rVW85XSaDexkPVrri5L2tJXHcIC+53gcwa//k8hQJlpzhT9H9ie6UMyjNR239WLC
ZF8zLYOVyoYo46TR3B4EB0L656R5i2fV1ZWfhPKYu1uvDLLCYXA6Bj3kV7F0T1nU
kS9RPnpeweTLfHSTPsJkqnfrGxtudw2FvYJ5mnop+w3njJp9i+2gl3Vig23+w0nc
gmqvjS/eY3WhxuisCsKPOv2TASKRY7ai/7w4O7MvjIX37zcxd9HMZHBOkdVhjYuE
5F5mwryfnJzIJ+3K5hU4R3gXBSygVyF3gl+VE67KEEz/zdHwttfaPdO0X4k1+VDP
YpO86a27aptGRJGUGbTl9lL5RcM+QbqNGj0uFto//tyyTM8jMms6jg8kVc2WBl0N
TcixqljvuTv1mr71KnHsT5CcgJO14C0YUkz2neXY5+mTtwD2p2blEfOasDtU23Jo
FHj7V8YTyVY7zpC/n4QzFbsbwGZLdI9hGiyuSOqstk3jQPvoSdpNQ3BVtLnXtmI3
OjHiTkNC0e0Sl8vhG9inKLdgvRFsSenCtBkDOKfhIVUekthd6hzRgbnlWyu4aoYH
9YOrC9dzKDiflan81XF2mBvKw4DonNJ7CMxA7T8mMKV6SSabFFDnTDgzM0Qw0eOF
vtraj2WX4rpX3QGF7ZNI43/aIJ3LSYMVfx0MiBcD6hii6h8HDhwrmpbgoeKaxtOL
Rey55bzfphzJEpzGyboOVdUFqaQMohJRWGKQm3SRYPN8sJDk2v1KOBz5y3t2/NYi
9ghfFyWa6+BwaD3kG9JDTz6K5xP48xJv64Vm6iUgQ0gTvhrXmvGK4gJK1+aMT2Ez
5P7vJrujxZpau610ruo4ZjlqKZLa+cGlJTqfaAk3icH4hoAAHrYksuxJyu1Wuaaj
M6W768OehF4bDH5BvianOEig5S5k7JseSu++gG383K5H0qlPU7m3euxLbSu2CNfW
SMuaR0+O7sYQzs9w/WNZ9JKC1ekbAn2wZtFMOhriA4ZUx67TtjyyquhtUcheblwC
512W32qQxTek9PMGW0POhomaoU9T+MyqhX2ageOTv0sejOZBTEop6GzbeoSYTzP7
yOeUgPr/C+EjxfOgziDuUBl1sMIFmjOBexVWuF80pqL0LCfwOPwkG8CsclhN4QLP
n77HOXAJjzTnR8qa2SZwcTeAB5P2S8/eJ8zlCYvUny0Me+If0ZA5DILr5yDCod7q
flsklpAu7FEAAMFo+BvRRp/b2K3YmktHE2cC+erDtI/hGIyvVEEp2OJOeeFw3UW4
lBWALZUOku9mXeD65Cb8yNDhLRZJr0xLu885afRY2DALWC4yStQigh9eBzSmtVL2
f5wpoN0WDvfPQOvCtlqAdd6/ScbtecaSf6HYpVwW21D5IyO7gcN31+Kno3IFuVuD
yZYi15NabczXo+jrfFZRfRRQs/X1FQhYg4APHzOimOU8MggZRnFny7X5ADr5DCU8
uldP1ZRKBZQNQbExrLUPZxWj6dPl+m7JolxGgFbplVK+aoNFYS2SRmR4pB6GpfNZ
nWitDCFDFpsbVkbb5JBe9Vlf88om0sszsOhtgyGzpE/wiIqHmud9k62d5nl+Ylx0
16/BjuMuhm9YHBmnMAdIR+U1SDFN/5U6AbStmTC6qLy2gaUY8POv3L6NKCwODWis
tmAs4actVCx7y5jNnKQyK8DMH8WNvQm4KieRanAB/0KTBlx4FKgSIZd1W8AOxaWe
U9Hk/UOQqzrOds1+0OSVJIT+dU7fOV0GKC5Ew8ORw5akPyol3DWUD7TXrxCREbNg
3bbozXC+Swnc3g+nsIAYkU8oLnFGF3V36s/iXnRt+qvO+02y18uVIQZ1gojPy22T
UragGPrhrp1T03d7F5VCGKK/abcVD+VjQ6Vt+pBbDMww8ZunhjvuNvNAyjbcI38h
9ZJUl7SVVNyJfn5bZy7YrPHShFdxMajRoh+c8OPuZXY7ineyPURSMFN3BHTe2FEw
1vh6dyRRggp90dmWU6e+zA+d0r/rtZD/vUMXDdA9F4QPrCSeqDEPY8DfGpjxCCVn
1Jvk+3K6ceX2BUNe6woy01mhVKCj9BgKuSjaE316TpoDPOs8zQ2nRKzTFkDfbaeZ
Rl8oBX1Bn/70xzLTQuf1xSAnH52nXFevC9AXCqwBt5SBHxP23IVxFIyi7vTEpIGm
nCgmuCRZbRqagAvaOwiozHDl4SMPdbQPJFdpLsB36uggHHIFx6QlPCjXfulOPljz
2WwA13OhW8XQRlUm2u7XYlSEuELJ4cMLO+70NnOigJXm4xgmX+2UP0jCsotkkDWX
pzIJ4gl1QUD9cLWvniyEXAOrzPvgrxxv/74hfu66IwmZhMCmjU9Vb8ak9GbWhl4R
y/0V4tuHRLDPnUO53bgfyRcP07pDTEyIDAHTiWYCxtCeL31fdjNeqT0MFEv4YaZf
mCUwA8kPP934cI2/Gobsc3DrLHRF2W9wgeQ5LzfHFvR21qF+Tiw0jLRgFeTWz7kt
MaodjB5N38N7HDPMt9NnoSEkxLby8MYz5c5xBp1jv2oZQIDJvBOuPdUrMu2vGXef
ZlrjJg7rzmFTwnG6ZgEOKVTLuguBOE/JCFaX3nJGvn9M6cd5GrxdT0Kxxoj2RMCU
vNlF6t8HYRW3kf379ZhWXCN4ihHZiK+2AEPjA6ThukUALZo/ODj1/F7iXMwAjrxx
3F70kearYG1/dw+22BfExVjkPrzTPtxV8P1JRsk90idypmalKyMZ7UHoZcPxgh58
7BDPL0i/WWUC97PmRCBFAoOdSVFg7AsabNjRTqHxalugfBQLMGbQ8n3D5h5pNLoW
yABKysDmaK6R5QrQ7VtoLsEJCfHs110i4mkPICOqDRMFb3wZUdPeGNGwaKearLBC
aoFKlhm4CrumLDDdswjr/3/tjQhi6bkjEz1GT45MDtZx20tKzAJ/uNX7DwNxfudc
v02lPLqdtZs2yrHPZ8ERwPDTPv0nfJC63GBLqGQ3NEtm9ItrXKbGSlqc9kJzDgyf
cX1nb5VBwbzcZhq++lAwH6z7HhM0JZHNm2KiOy35BW+0XyppZtxrJ1GY+ut1jgZS
33CsixarZSLGhmoxiMLJ7FN7tbng3MYTLun8UX1k1IN+FFVAPhbuegVZqoPBFaS0
SVBXS6f0/yZLrRP2/2Y1zwtkRLfsItJiV/l7fMLpUFH/Kcoo4bOdpYIfXl/bw5uX
jci8cjvulCrSP6a9Qt8iDzG4Lo1dg9wnUoTH0FaOoCG3IpB4PD8osMjftcNUDfXK
UvBxSsoU7+VOYTUESYTBItyM/KZWFR0oksqBOAxXoFjbIIXnhVCeQOlrcfEWX/Wf
pF3wANnvs1ClSWzIDNRmGAK8IoaXoKGBNeElpZq617u+DkVNsSR1N1p8ETqSSRvA
D8FUf/bF/z0Qg6UuOhIl+c8n9cfoR5s/WY43W6dg1I3l2ZJMN0DVckqpa6BCCVJA
PxaiE5Ul4IyPX0PrEzdu6Q6jffTsooO2F4iuduSoL3/9LirUlKUirHyrAd4EOs5A
oZHftwQ/FwCBSg7j79T2EVwPpz6+/vdo7yymdprZCyzbCpTR+XCBhtguIXPhmxD5
Ow0SXwt0j4C4eXYqKD8gx7yVfw5oPBneJq4grpbTqhBqaOq/n5m9kctEq5FDBGvc
pz9OgdvdY6+cKt/6GUkSzNVtlhXCGQUcnhJbUajGPqC/a8DQyif8fgz7WxWclSr8
tUVxT9zUWG2MEaABHHLbj/u6/dOe1I7aosil3u1XbGD66pN9v5+ZSLtpodBno923
NSZvHYjHbML1K1/EojQmISESgfgz0zIOFFH/BeKzHUgT3cjAhp2SwLcN1+pNvgEi
U/NXYMno2EqhVZm2MQi7p3DN8OEpt2Mgn+81UjZDYKZTf+Rt2nX6jpmhClOs1Ldg
SmO0oORmxC6DtXyk6x3P0Nc36Nh9DEwc+029As+UliqD+SX/X8yKQCCfL0mhOfEa
DTsrMd+wxOyPIT2pLd4Qw+hwkd9nSsWZBSD8WSstyZEv7vCCV3um+XuaFkAHHBnf
mQW0nisQHALJvhLX6Yz1KWLiiC7Zq6hDWBY3yWU0XOLTgz60gMVKsQej7JeeX/xo
+ADHq36h+5zSo/S4PDXySDUu4XiOFZ/WQpKd6Akuf4FzKVIDOdaDo4Zac1Dyoi0A
OpNYbmR8HmKCxEMs2cdkTDVAAiJt9p286tJsWElQ6FwYYKWAc5muOrf+FYjP2xha
NYqjmn12qb9FKViJDjVFMTZh83BhWCs0sGd+yIF4QrBztCn5d6V07Dj+wzYbzpR4
0lbXH5R7E2dGT6dxHfw9cM8G2ZgrvaCM41NMkLdHMYoHu5RQqmXeuE/84jQ6V2pb
6JbRvdagQEf9VPL+YZ2394F+32EuC8gBGgRZG9uwAz7WczNtJ/Xbrnd+AA/nO4oi
4XexfwVN8OCdr3+gsEwUwl143vms6It3IKTgcYqhOyVLG3l9jloS8k/nPMVSqNSz
W5QVUQYbde0qy9sJh7QRuw2sPNmFpPrDyL72wCdvjwA7GWnbQ54XcMa3anIt7Mov
sifv7Becnqo158sftfXxSs+ukl8ujp/8ca36pFgv94XTZFRxzSOBv0LgYVnUzhbQ
XjXGshUYbORP4db205wUd5s+Gv5rXezDjxfts2+3jwOK6sUnIzWzJnORzyJdStFS
kyBy92ThAhi2JqMlQ//P9nRuZ0ZCZyhSZcusO0OuwfWcsSjKdzJZeyr705p/pHhb
u/mtdgcnwOE6FyEPOnrqnFQK0EizasoBPsKm/BU0CuunwDN3FidBLB+z74WwWaPI
+lne/pFQqIo7jVpNYgYRT3qXZEj8S+AzQYUBzPNc973IN2ZZVFtCC22uBtdTJ5KW
E8v1uqtn2JmhoZNAjs5p5L7aQiIpOjWNeVq4HADNwSZR8yx63qJDbT3KXpYs1bTF
CcFudYsd71/8UhCADv4DtIBtg/FD8YfSG4av9p/3LJF8fsHnANx3c2GBZKWN2U5U
JB7C41l2Xg9vH12hkX43zmpbMSghrjN7mmPX9j2Wy68wQfjp8hIpw9PTSF/a0smR
ZV+vJpbvBZQoV5kA81p4L7PHhYtqYV+Z8HAQBWdI6CGfdhsLHZYXJVt9c3p1YmQ4
jxe1r0u65/5LImTrjAUnSAUsKahWImB43cgvjFdf/dVW/bR4ogSkFuy/K48VLK92
eyNZnRtyBppdofl8Aj7emFGeYaRq0gJO/oGUigX3NfGpPK/6lf9QlU14T5p9mxYu
fbNEWx9qKHjDfzhjis1sAonmdZWsdpEt8Pmsw7kG9J34i/yXEoqg+kme8UD4ppJN
IFuwxRsIwo0HAcJDOJm8EmG6vAo6qiMLnJGFdRLt7dReuNfZgB8xFni7zk4o/L/V
BfzNNZYr9G/6aBG1Po7WqQKo4NysCVb1Xl5lQHFG3LUp3GntaPYywxRZnIVZoayc
TdCaZ+7rS3XxSH1cum7HGBEi8a+S6n1iFgyaOCSkkNOa0uBLgMRpGCJhx/WuNhBK
5kRFLGeci3B7u0bQ9iu5V8ItQS4vli+Ue/v9ftQviKv8lLMUJbafRsvAPrMlHJDz
ea2aK0jHP712qNjFUdIf/LESeSuP5ptlWI9Nm/5pOuHRx8GbFeyWL5Y42gJcBtRV
CySQJ+AQ2gKkLQh+Ds66QJGX8gIF5FVHitEe1BA55QeqH8mCBEJBvhNxCNaDwo4K
x6N4evMuxCkOlI4X24ThXvkSqMQRACLH0w91HPgIwcbjsVVCE0eNUAXCazuBHyO5
dWPcrKQzGAHGRdHSdB+qNOZDS1r3q63UmRqYFmmyBpHCLE5PjrpH6hkKd4LOl7vL
k3ajOigkvDVRBq1i2tqF3ptp5bmd8Qogdo9RK7lplrSKyHoGAtl64fyp9b00vH5I
VFI7+PMefdk4k9NtbEg1fQClhKOeKdgiOyMbq8+h8KPXWvl8I811LYv8SQkcxBiB
4djFZ0x2+QRm8SjOOllpoRd4umjM2ielTA9xuusucH2gjUKy/slA3k9OjQS4whBn
bS+Y6EXDOURGTgXxbbbaGoJS7JxMh5xE4NhBjuxeVfWuBDDiZwFOOpw5OLIsLuEj
zs7iEgffIwxS0e6Yl7s1fJd7L+CtpIVxxLJTzapEKZijnACYsmXmSo3/i/THSh70
Tty1I8E/hNMmFs7z7Nh57sKTGO/7wSjBcBKScpbtMXg8MCHMj39lZsBnsR6yLiho
aQkV9EazV0bphUooeu/qdztUngf6t3ndqy/TYhm44Id4ga92o2fyNoCB8aB6ZRkh
5douSvhD5rXLKj2C7XPOwtEBX7I40S/tjCljHBcwV0v+6oeo9VnkBaL04G3OAogk
fuiGRUOuMkVivmeT78/fYUWKDISC8M6FHHC/G20pQmTou5dIdJk9FpWM8U5VOs05
4pGslB6ig62KAgqdrXC/apzwso8cXdJbdC/9Wz7bKfqnee/XaPeZtk7x2YlWUBUq
d6GFtBveQTHL2SRZi4bLPlFeFRyaL5wJcLvFxQiZgMmTnpSw1w5cwboZ3Oumn2kS
/5qfa0hwmUR3nSRy7wUXEAxBVrOPdvLMYnbcPSI2hswFbzRW0yQd+XEA6wrEnv7m
p03cFgXXEHVoKJhTixin/nPYtaSFeTC+raVNZx6MHZaxSJ28xU7lpqiNPVzU7Pnh
MhPdPShg5xE+Wx+IECDQ5kVn+03m/CTRY6l+8gqWC8avnIAEDCQZmu3LvXf7rjMn
iUbe0YbCzM9Tg5OsqzUyozHQbyJT7mVKXt94CF4Eh8dCi4BbXwA0GJ2sOKqjQ4Pb
xc6bzFSsaW5QfFz6huwQ7OHgx0g4wnYuftGBeZRflZ5TeH7FLpHU2xsJQ1ATf0u4
PNGuvHoez+jYpn2wBS1DKr7rILifvqD+/6uzS+wN/a0JoqT4ALkr9o8h/PElkAa6
u42xpM/GtEKhQiNlDFGUD3+tXt479hHDkXgrn9osoj+Xu+TKlJccv829ilTtyP/c
k4K3UV6MW0aTJCLsPwS+P/WHy/qievfIbh9g3GyASXz1ZOwNy5XV9yv1WtlTuLUn
S7TRmkAmV5z08rbh1rJlbkmtB+rMdAf1KUyOrJvI0tXAumGoOv2MiqEEcx1hcPOa
zhd2myCn2QuxuL0iiUalUEo/q+t+8ZVDAqC+MViof/c2BgQTlvJjJnTrAGwlI4Rt
jTT8Y6TaMYutRUPfFe4NrkQhtonnd+CI9TCYuXb3KUP4zZ4EvipsZj6Uve4/Mfoe
c/JJxCBMlIP6G55ZvWd0Tjls304u5ipy38qmHpU7LSvImol5hC6uhP4EYphvf1iz
OIT3nArmyu/Vx9LK9LtPK6zWF5LsT/GH776gYzLQ0hszOFhcLhPAi5hvM4KV/EMT
JW9PrMdmVrXLG21p+fDBy5i+mU/kgJUtcUz/aDz+H/ENTQd5GkLKZ5qKkkYdrekU
tndQVk5PdMSgK9sCLRW0wQznS7vCzcFfFMIzwVepE090ZMyGVl63FtFc2fVoepBd
S+f0Vpdp8GlxjFGsZQ7ziClJLIcWy0+b3b2SEQab7RXr0y/Th66S4woKEe+ToE/u
2lc3Bd1OYaHO/NEaWp98Bg9ZVyn1IO62XimA4I7BHtpSIWUDYTLnrG8eh36nqdcR
XATv+7agOrPiageynJw9Yzlicll+krvCVkQZ7qN/y9HpH7aYA0NCzOrlTGLkaDh0
Uqkdggj3nMrzAOPt8pvqR+xJBCnvQI70NJlsV9xFCDq9i5jYA6h4GNevJMVBg7U6
Eol10xfDm1axYGsa5FRupIysDe6UtqegNdYhf1mHfrLRH6hahYTDadcgKTHwXPAq
6ht1teAOCNeq1sVrkopgMzzDv16u8POOPH2VbPKAB5e5LsPxdbVi9/Uv60Or1vat
Oo+P755OdynV+HmsOP5rWUpNgMjBKPgRDw9HKYBn7fpVAR3PayHyoCzKBbZps0P8
dILb/0WIDiak/5he825p1EoJd23icu8XCFckdHzIkyMR2KY07zbXy9y9aUWnSLvf
3HHkq+QEqpZtO71RFHgaqC6+2oKDU4cZtcVCnxJWK54lZXrydsjYOfFLuOZxbaZ5
Y+cP4HxNb+zNpR1l/FX1R/+J/h0eeaOpkV7QWK++jf3St7+zGnEePwS7A9Loqxxf
XJDn3XX3WfVMGynfT3HX4aJzn3vha0zbMsrfR/VzxhPAlFu0/Mo9hDt8hsjOcvoR
4nPHLC2q6AT/Hl3yet3h4XdzXvJBKj37qFD+yi6bBIbqj9bSzVQ0Z8KuVcVwP9sH
rNZ19Y5SLEr8OdNNe9JvaZ9DzwutRt450I00V1mXIupXO8YOJb+moByPiRKwmP/h
yMIIpRmPb/wXqDUbtzOj34lqXNXYhBF/2BjXIJxw01BCaWYke0HX+6GECXLrlFOj
eS0/TAEBSHterfsPQVWSlm60U2kS/Utuvp3IZ4heagzkhUleiz70JSrevnI/eCbW
pSsENGL8niBaq5Ib3jsMIMOMHv/3ynj1r+PjyFCLKgQ9L5uPJlOV3w/R31D3JWfr
X6MzkyU7odqhANBetrDiP/DURUqJ/z4AEIh1kZsiB1cQ8UcP1BYqj8uOqUMCVgfz
9MdVwGlIcO8TlcItplHsBZ0QiALP9koTA+WfPI6+ENWvemURHxHPmUGAtv6WIwIC
zsUHSdEbRPJbDg5lLUTOLsCxB4NZspKiQt2kHwOdMZug8L5jj1DKBWc+CpjE0BJC
eyuUPcuMZMiOgYyYLfLirepIpxH+8BZkl2a/VQoltP//Z19KeShNSS6ICotsXUWb
3Af6RKVcF52/pMjrHWtAnYW919hW1WQ9DlUPX8aJ3/gBuxrd4OigxRm0ML8Z+4CA
1T5g8Glgy9HMzlG+8itVaMAzVbEHcCN66DnP3CTGfmrpWx+kiD2O7t4jOaaiVF4W
YA9drlWtIpPjlNe4dMWhuQ1qfw7oOmKhBG4ciem7lqtP2wZf7eRDYDkAXeL6vA6c
VrP7W/nmzMCJdhvucMlxDDLgqxlFMv9dHXZMS/1jKYwDjyON2+d/UO/SjpoCoFUh
mZIhBp1Q3TWgfgbo5um/ZD/FIsYJvdexJiP421jauE6J5PSouUfxqWNQO3YN5qIt
hZFOIUCLfrvy45ErOXYbccJx9PkRytUOmlh9hX9pfayGr8tLa/l4APqFZqts3HoX
LfBnlYrqlfdpjdEq+2pENH1m6KBPvOn9fOVoKZJxHeATB7ZAIaZKhjc1+FDTp6zc
zKUSwOjDK65k5fsjteXIwVLdpNUt3btv+gcJUUIndwmCNo+JKHC1UcsXDRswaQhT
tjqR7cjibY/YuZiHBdGVf8KSBXzLDK5i21ej/4aMps2n2Fqec2LpWU/0MyYi+h9u
ZXuJBD6SrdxGobWdZ+uQ+1g8ko6Uzrw5k00rbY3K0qfnfgqndDEXmfVLSPYs3pFB
qsDH/qmbhlDtb8b8OPxCcLJqCpYLBjcTleTzsSD2mmlhZjkTHrWHjLQIgvz6FQLC
fXw3oCD6Paj4/G7WE6fp1puFS3Ye/bWO2DhBHArYVaAKi5zJyawAxzgS1x37TAoK
d9vxb7RY8nzvZHPLxBsN6AXQPA9syuK+hQi0KyPKhgNQ/GXW3nbuPGDzWykCkMTX
4oMFqYdgW3oXU1FXTlrDjjF4yTvbU8y+9lywGYHqDvJuFiLpfDzpyKHBaxCq1OeH
nGymW2suX/zFlwf17bP+ZB9g9Vk5hL3VsVP6osZiEKQvJ//Soc4LCzOR8AFAPMKo
cJch0WGj216cm1H55D6V5hcZ1PI2n3F1tnU0F88iG2jWu0a5PUYVZeySgy9+gpTo
VZS8KHdEMW1TW4GQYEGFQZs7/rF+WbI80ToCxFDfJBzYrcTKb9XppRjYN45A2NpW
kYU/12zOJv+BwJ34L8WHMl/O8o24v8fqNqmIkhOv+BkxdApC6BGBZRjPbas/5iiO
2Bk/JVkqeVqGTvZ31N/RtUkG152NYwnfxxTr1wcpDSRVvYeEpt0pZzFiFjzaj6p5
ucx5zC69B/FrpJScUzBoszf47W+ZkfVvIlj1ZXQrJ0KHbVMJQBKg35NDIZEXCwbf
MgBuiS/yPeo7RtgNyAIRG5boXsjpUpXmsH6iMw3FpuTkjlHNmrvk2BRBzyNTDbw9
pUboVUviOrdqKflYKvYOTiu6fswDkP6wCJLhlaHD463hD0Rf+qQpgiJsyLBf4Jaq
QEUAnwjjxB6XbK/oyY4m20/QgaobiKzBn/fEG703LBm/WoMvMRNvGPtt5Kj6Enzy
DWvcxeaHX4ueYS36nzZShkSy4A/zTtL9Kb9H4Fk/1UGJJloRfHRUCbUi8HIJ7AFZ
ZbODQu20Z092OHY9YHH2IZZp6ypwHqzgz/KWBK43Cdoyxp0eduL+xy1NZdoizIZm
N9JI3iy5Jk4oT7VMkuic5Dmk43T7Z3jmOIvyOM9CCyUwzU3Di3ElfRF58AEahgNi
AhsrJOhcWNeNRQmcayhYtwOZrK3tOeWV0jyemGPrRjs2Ka8ydDRzkMMU10IGUhfm
MYzGZyCUl1VVS+4CGlRcOTUX6KUtle/N9I4pkI6d4mcRqf17V7JGtqLmzRS8zxw3
xnykqo9xbe2udyV8yLj1Bqdr3Ro3RbTrdyZzDHJErIszInUYx6mNIW0sScQya3uG
6YzyGIK+3eQeCBkDCAAahBNryiEEcRKg88Hi/WHtqewPI+4rBjqjcql2VFP/rWhl
ww0j83+e32lhMnlGDtuccsNy7ikR8rSGzrvLV4/YjAFq9FmUS8JG8AweYKeKC9Kw
BhZrGbLNb6inUKm8mNqdvLBRRlcQC9vWMG4DFaETcs9ctrQ+02JLPIqiQdUxudsD
YMZN/Le3b+MKAu3hviFZO3YwRF03XL8RiPmQRYrfmp3Dw0bF4ukSli3Q7bWAAyNy
ONsKt80SyUuPL4PtTC7x6I2cgdrswQl6jjtTUIC5HpB0FmQres1kW3PB5olDyuV9
k6F0y5jnCBSeEw5I30GnC2idVh4aWbjZHLzwzC0fqnv1lPeXQostZUJx0AvJ1kw2
bPiV9DWvZbD2LEzlqWAorDSq2ebKFJHtElaQlert2i/6D/7IYTS35IVqubZ7hWr1
/ZWwkUijxPTWg83mMUP+MlcSiO+RUGEdBVsqh1ydmPfyqMBbDMwPaao0AaYdN4QM
AiRnZP7mEbOsPl7snEd5RHMLW97ukyfzzv0sPBdjhevgzwTdPHC4htRMbK7UnR38
v0rJ22Cq5eiCHynFbASaV2LB79inrcQBHmUUKoOzEf8NVsiEBYs6Ngkkf6zO642o
o0faNb/D/3w4y7ltbgo4Hzv2Fo0gB1sJUEYKrwNP4XDsGr6sN77aeAnrQXzzvqKP
Z+NVFx/yjO1KtE6fksRSlITSgY/GyW/iRGayxnW1rzptJxohPxvFqksRyuA872hP
cF7cKBbS+Y82bCJtJGZof4CZ7W2hXi82C3eDjPx8koOb4FBOti/UxsyPwh1ILMNI
PHoU1gPLkzXP0+K4tgQaHHi5IrCTmFTOPl1/dlDBCAQ0vFdgzJucFeb9QTmIuer5
JLyd8sMox5pdtMTifwNN68VfONy05yHLRzlkJqynEoJI6XAHH3dywZZOqbrscOnP
U181DpYA5IXgPrePlpPVwTVNPzhy6Oeyfm3U3EPmdYAjPrpqJz9TYQ6/P9GozdVv
9WezWKytgxFJ/Yprp0DiikmkvC7CCFj/zkqnaZfxEG7bYv/rxsdIWokKjokVxHO6
Rm9xX31NC255tfQK+sDRfv1WIaxuFnREqrgvEdOAbX7Ps6j303PcyI6ZbhUuEWjW
Fth/ltjRBxyLdqzwPyy1Dp6C7zTDFl3OOwIOcx+qKMfeSXkW4+tI7oOGvI+DkBt8
+0C1xQC7KzBHvUc2a6CbEj41QkjwAg5bp75H7raNnaN3rnbAm0lehEuCsyMLb61t
KdgGoAuqWEHSvQuU2E7V2rJ6APPEzsO67k1ckqDT/2162MLPz4QR0JaMOpw1LruL
htp4iL4/zZB0F4s5iqIsxcgKJDQHOdXY7oOw7YRO76yfXNNN7YSUNCG/rS1qn6sJ
p9WArYtC7F+MJyetrla9IpwJpPHgU/UU4M2put2jFDAUrLFxvIHZUzwornQMm8VG
JA4OF4Nx0BmqETkzmYoPD4A9k3QbLmyj+18XNqn0bZHcXxVzSkvV4pF2lasMrlgx
f65HyLbcoG2smTwnpEkMqpoWTzs3aqQnN5ogxSCHm3Bu8bJN63GIQ0p+CWp+Dzlp
emcPAlZ5P7JIo1JrOMFaowoQqHPyQB5gD4UFpABif7yMHYSuymKdZIinMYpP9hSV
FT6WERSE9iTzoMNP/gVxtnvsUziAgnvgqFePzjGAIZCPR6w4+qI93JlF+iuKjAR/
uDvXh6SVlP1b/GQVCjE9my3YbALM82pQd7mc6qZiArH0ipRu3/oFZUYKDv9xtlqf
V8nCZg8WgzZORiU4WAUCxG8+ajGcuMHP397U3iUpID78qtOtRdy01mDafqRzCa7x
LLG8fR9eLq8BhVKQGvHPZ/oS7QBRh/RHCkAHncEWjoXdPg8YygESZJdjfzHfxOS/
hWsIBieT/QRvUdVr60kagoBYK468BhRe8M0xt4wPFzbGwosxXFi+zrZtz/8TxF34
ZADaqwLSCO2f8h2uVdr1vSicVasb2w6fBzqqn1epjHlqsDKXdoQEvujgjEdMmmHy
8HhWxj6b0DBD7cQ/x9pk5aPmlldIxqhGoRxWWcsQRh8iWtEV11YmfiMl+rpm/V2x
TBezpmwf0P9y7ZoVZYMuMPHWwwV0ECQIKEq5Z76pnGk1V973HJ3ODH4dGD0MAyus
AMt5L50xY4CUvqyT2WNfGYsX5oFUw4aBtJsjBoRUrvkAixfgAgRz+TTwKwhchiUA
glBKWIRFo3Rw1fGwDhNk1qxCkiDj7IQG7iwaElr3KQ5EXg6bqH0air/b7mUhk9vP
6RCg5T/I3oaX8400g4ACmd4vRrWvLUlDsaP7kD38UUg789qzCuxtDklR8S9qI6Am
vaTJMMyQXueC3gnG0fH9US/0zoFni98SUXx9rvuz/s2tRQAaN83uvR8qnjV99AaT
WXV9aPH0qDN491A4AG9X2yBh27wG2EdkCPTmTktv0HAmU2c0Ysx6elT7i8y9lrv2
ZG1RBZh61iwUpiz1SEoOJtFrNCHOYy7u+0XHKTp0x93puylJXNSdhtST4FKdoxel
VvHnSEfjGvZV3emmkv/F9aaaLm/RNqfn5vgqB0w+XuAobxEH98E+xZyMzvfUWzdv
527Lz24dnM7mD58Y3D4s+JkvMvPLNQijRDkAcqtzMk9E6uNOXFLk9Guci6jNnCIx
eqpmq4o42SXataUCukAujoRSxm9iOFfzcsPTY002xGCW2cDm4nMJ5opWNZ7rvJRZ
edr2J9U/b1gAhtQBPv+Cg15af7dy+mwit+pOGZ1nkVWxjkx71Oz8tnV5X+x86z67
NxnVS6bLrG9S7NLbFG/nTsOX74JTr5ihJeYVbZnSvvObaYUxwZaq4LgNRyBhJ1Vq
qVj7gSttNlpQhPqtak+bSKy+aDxHiwKbOzYLJx4d89e+Kco3jRq7P7AXfhl9XHwS
PzqRysuCOQgmk2Zv0ng1B1w8hrkowIGZ7HMisvulvSRy2VkaSHkQYQAPKb06GsU3
aIPD4QUm+7C5dxmBvjX2OtOwoPO/MXQkztRpr0UfgZ/cNPTlR/BA8Y/Ck9tJnv/6
QLOa+2b9s6s2QzVRpZzJC2fMjN/7/ekmazKeYtxiT5aYl7zKvYLfYlv1bzlveTi1
21npWRD/VjZiBYv4lwwUodF84fWGLPU/IJ71PvkquyqIMRXYkgcfcn+ijcb1ABl7
G53x8ULyonS8Q74QyNjqSnYaW2rMHYu8/zSQxb/vm/FUQtzxYV99dw5XvAdcDrnu
c+rqXNmpDfQLx5efLj7MpyDTHACjrUrwTGs0JUt3NSbwlctvidpSnl8eqOK4iixP
6j/laJlqddQBLaJm75rxMZ9+67e+XqSCfimLxDIXd5EO07J4f6rffCDdDrNokqqR
Cj685/PEg2GJtRHox6rE5GJ0HzxHCWEHnc1HM3dmQjDpN1ItLgk+ip8d5J8xVpID
el9F/U+1eDFbxk79CPvQBbXqKfvhuMZt73TXB5Wet4NGr60UmcZO45QIiQjzLBBG
wCnjvRYan5aK9nPraPwvVcCweo6UTscKj7QisBDSD9asecmyyfMaN/8Pjt5eGCbY
8X5ry+IjGEzeWsB4c2iJwj9YXRw7btoq+nlrzyfky0HpoIOA1Kkk+9tpnarVzpKK
Nk4RaEkqOTSdsEI28oRrIRbendGPRsoV62X4rn6f4Jx8fivlA1+zNRvF30IG7KD4
zWqp4A3/p92Fvl2fY8F3B3h9qheIRN0JEAsXGJrcTPJTXHEyN51XdmTSbzu7F8AR
6b5Vw3niuvekL/sHUm/nNT9Y6Abn3HOedqP4bT1C/dIUxWlEr9QSG+R8P/BlzbmC
uzkZ+EsR2pOslQI6OXNcmErLY+RH6vbko4qRRhGwmvjrBUjDGqXMFpMsc6z410r6
cxx9CMpfq2SBDSHFoidqvVDZvDz30JINGxi03WOX+vqPNqwi6Ur8V5TDnUIo2vqy
1feBYWYpIM9+4u3Y6BPOhqFD9n83NgeTt5CD0KXeMsBwa+1xenzW4gyn7hDmYnGB
hbFHivh4Nq0pKWlC8BKmQ7OiA5XSgdFHKoHjV7plCdhEfUg5KzmLnq/V+jKn3hlr
3YT6j4VSkNtZqWwtjeULLMgLw0SWO1HXYwVCkdOPOJfvvQMotdryBFE/2OHiaTyv
VY3emUq38X4//d6ABvec+ecznkQTCek9OeSaOg+0OP8z2IYYJ4KGwmNjIX5L3x1R
nKluLx1vj6XU/kAveav4AX3HUjGDXXyp19z/4YipOL1lDq+ynN8mHB2bFrZ5rjO/
RtaM9iP/hg3YRaeW7R983lXryE1O63QxaP0APFZ0dmWqQ2UriS6kSKCkJhZIC5+g
m5IJc2scyVAx7uVwkLwhTEYZoXWfmiftLqcmBOhviyfXXZJMiGlL38RWi+gZY/qw
QB1Ftj7FoGbDczJ0HsJM/doT97/pc0ajLDJtlfsxmLPjOR3DT57usFIaLh+OcSUL
cWcMo+QYM3WlV7AC9ezWNpv+CfxQE0GXxsYXp8WPSBYR3gg4GcGXbGAWYekb5NdO
Q9aWMhE08lAKOE+mynZRzaNZQKSXJ0hLfI0ygrIoNWkiw/1WoIffU1tCdzJRajzf
Y6LCQr8jbN2JeQnGJUrc6o3g3GPATNXuV2y4eu9wWeyJiFM/rX2RQu5WLA2/IqGZ
JcVE1HsMuFuYc0X9P+6bEqTgW4mJoTcyHzMNEdfaeChk6AXAIOl5NrtjMZxlS5Cp
MvU2d/Y3NlmTkBvhnnDsHCcJx/I8CpArJREDYBg+Ena6BfNvvmDMierUcCFsGOHs
jvZQFk9wSs5OlXin+NwMYCLh6wa0sP6k6W/NmEdGGb6mH/MvEuqY/MAzQE3nwG44
bMtMM6t6IXGkV+teQ4B8FIRxuE9eXYzMo34+CTI8PrRrq4tzPu9c34sblmvb0N4D
0EKrCkG5jvcyBYze/hlCCRSzV0tTqwVCmlQ9lFJj4kBS9JeljanBSTxa8mPcIxdf
JwVCH1IVfWtquw2KiUtZWjlCl+lDrJVrn3DYMf0vAAq19pxwtDnVN/yfXU57l0yJ
7traFyJhiuZLVGqxm332oMsP1ksFz6yqmnExdp5Hmmb/Qwk6/PQFzXNnyMhkKGYO
a0qPxGUsUeWDdNOecpQeY3gobSkxua2LzMQRLbZamaiS8/5SnhgzYm/ncQYj6rYg
/zFey73JJJoMHEOG0kIgCIBy7CxLEDP6XlyxiPt+8nnZiyfPFb5FXdgkJSjNgUQc
RxMBas1e7tQa037SLwg63OmXZF0NJ15wHnu/vvRfktzRsKVpToX7zdwnJpcU79Tr
8vfkECjvMy5L0oouNTdXy7u7wp+gui08gfYnvrucLDGYJ3ZgZxc6+M4NOLbYgJun
MAQgrugbNoQe3I6J2C5wvtDyhoWjLZPd0O+QbfJdNt6eypBR01AOABRkBtrvuj6h
uPAkhSTMSozVKpVHt+1JDv7zUjjAct8jdLDWv460VC7IDTYdS/RKxSfi9Gk3ZPY1
wopV0+SBT3jsQa9cdgQb08Ogv106mjthdIL/d1WZiUAjd8Mzv48sBFNvD1X5mwNe
1o77skvutRItGnOU6aSGtSDbvCFV5B6J4ViEF7zK5M8RcoY7iPEL2ZHskNRliX1o
4kpFF6r4bfVt4m7hjdYz3mT24pBrif4BOEF6rNXdr/4c34XHifN4+KRndmn7lPIh
wVX1fXwqHF1+25jN0cdOyfSoe4A3tQMG52/Fnld/NuInG/Igi6vsdADI7PEDJ0GX
Ar9IicyGKT8G/hk4h7oYC4mjGZbEMq/6lltIilCX96UOi7r1597X6q6J6z06IE8z
xUWwmMi9VmRzYqdHTSdnGi6VhWBOPAcS5iNWJHkV1zSc7bPVJJdgJkGHQ0SwTZgZ
iwxYRR+VRAui7FkqNh5Ou7woUKY7oNE0Hr3gaZam8utQYndbW+okIeQ42hmGleMt
OJhsoe/YZGrmKJ9LCRf0j034jAK/Buqa6PmEmi72MGu5oURVn9jUWUGcNam32nMj
GXCe0spKHdvk27vI7peiJLNpTW/Qiq+JsHzZb09DAjpewRhZARYHhYW7xvF+SZiv
aR/0dGZsk2Hl4LLwYWf7jFAxUctULKgghXwC5Fq4JcJbZM026ZyLuEygnaNgfsQn
B5JoQ6XhNh3Y0clKrIMFBO4ip1LULrDtncJ7c8vNa8dN2bxH7mE/9mnu9wTxStxE
LxUmRd+5G1P6WpD1nj8UNhdQPrsULikTnMfSc1COTu7N5pgTJdl3JRzAztap93Z4
kWlLCJ9omzxeWfq1TFmB4uGpRId6/NuMf4YnOH0HzYgTcUjz65ok4UxhNGg/u6LQ
7FsGEuvjPZsBJh5jfJYuVCgWIP7UYV43JnRIIxUkV5u+5x6sCqNuDfhxppD9Av8b
VuaXh29Qck/ULGaRc2kSwQPq7e3fM5nzUl4p77vdPnY31SCF3+gIggju0cQft+Ua
E4+VE5xIYhQ1VMsMLVMKd+woKKl7fcUgWaOfixduUyNS3GFU0ZNOipRK33pUONNi
9WAYoFjswZC4UUzyLGaaPSSGdQdCXjILnSIWcZUVZUKGxHyRM4rQao+aMUhKHmQb
MrIxJ8uq7VL17o8wz70THfaPAlozO+atP+0MHUgB0cljxfaKLtYMC0ynvPpYXrMh
xTXT6TBOJJa3WAViM+aPEA12gRiV6uqDICmO+1t2NNia5YaQ/MfMGHA4MUnFVK5t
ezrzsBf9ovGbR5zY0fIDjZypfDpCnuhAYQwXFBZLHLAaMVVN0iEaES7q8IDni8r+
y46U0wgMAssvbxpGfqobzLQPc0hFutgjRIBo3CV97FI+zGSZEJoqj9nB039XEs6C
xipZQNp7wbfsrSMmh9G+k65PGUnTRce7vSjK0DU3FdThH2XjL2HkAs3UrmKI1TfD
C3HuyOsgRtavn5KS/okfmK8rKE4rL1GSt34XIuQLWro63zWM53mp4XK6C537s1m+
tA2skluRUJTYW6TuwoTmm7/EeMwCN+Evv4zIwd38SAb8fjsyNHyxkiztXhkOEhfX
4dzzwC+GhqLcJ2V2QzO1f30MMwuzPFYK9xmCgmUmQARq+WQJVHl7So1fy/Ud6+mW
ZCSCtxw9tgxEJwAkQDYJNsNJ0BiMzsZtvNk9/Wux9+0XEOO9TkE1YqBASSiLCj7j
67XKmzNzlLF6LTWjV5DNFSbF4Uatv+kzW+C6XP6PoqPkd8ZEHScV/jzb+ySen39O
23qTufNkb6SNQJECNexFWB8UDTdvaDe6OjwIjijxqIQIlj8/3tduYKRetJgq2W5q
NTy3vScojAqGOIBA885jqGqxwaWggkaKfHXEJqQcAEz1Zh45DsY2j534+fw1x2cx
kr2JPSOISoT3+/6mCfyaNhGRaAOBES7+k9O6uU+km0mcWwaWEqm+QMLKbR7B6gGW
fQw0bifqO0BGBcY9ImKRpC5kfCYmQx4c0emUpgJwE58W0pDV6nZjeUTIfF/sKl8S
LOfrDLDp1b2F5NPy1879UDPwUtBAlTPs/5Zb8HIC9cUsQkjDrgph+vdWnxboq6K/
7T5t0h8lfxpYEDTWjVjvQczNzuPFaXNl8woxYWB3PODZcZbrwTcktPtzdaRcUKht
SE1BCWs1/OiC/5jaPq0yJO0b9YltD5mWMDavMbMSk3GZlKH8GPLzKwvnutHcRpzR
+Lvfg1V6RJgQJc90c3B/T0h7Vo9PczemrStCYvvZW4vcMost3eqnGD16KTTbbTT4
aOheaQLJUYFUZ0wjWzzFpVevtj89iSALdhrzSwoIUfMssweTSUnaslSItyZ0k4lF
fnGpucJ+xKnwHBxqxmG6guaVegKeIBhIssQ9ipHA1j6xOfmdEiBTbU18qxYSSKIn
jbKz1Ga2gid+NlYNxSKIdkGNNACDYUrPUXeFHx/WdzVApAdvSQe5pNcM6LeyVJMA
YDQsmBGLxNlNc5klYJNVRuHsCLuaQmwOmQdMTKSiTpl/A2ulzvNXrTSUY+8pxCR6
5AIC2Xp4SLqleZ/zWP5Vk0uHAU3IgjTEuknEHWuUQfIWXTklYQDB+5uwO+bdDU9m
SqD7zkM391nKB3roApHMwRYaNC+WbyMW+j0PC72RxxhvMqGiESBIdG82C2TOov/J
ysT0QTRUjvaUNPWEsSvLiqJU/kji95/ByF1+vKTXvUXlWDvcDeVEH7H00ptK6k45
wmNLFnoM0p/Zt9Vzfjb135fIhyKoOO/20ktSo6RJGCQXvHLQe39/uXc4mooKwtli
t4a/pp4W/BWDQ+ZKM8dDkAFTvabZzrwYMgR7gTsKn07Ku7eSKD9e3bNc1qS7JhZ/
OnNH0cWAjZdimZJ5lgp71uWrozT78jcm9Wl0FA7pIZ8qGu1LQXhEQuP4ROs01kJo
UTWRFb6Oh0KNd8aS8ghsklgBvz7p9usgR6fsFqJCnYWy33qXVfSUYz/BQRDKKAFu
CxUpEhh+CgZ9IOPUSkfCo6TK6j7L8Jls1Mug6K+tnftuG+Fc5MXSjTYD/NnFKPUs
8LKh1LUsPFENt6ibx0THZJ2NeHJDD51+UoQm21Rp+3dBmU8KJdY2v9z+UJvHLvNW
Fkz82zlCNiqkPH3hlSHfHeFija3KsW+cWgLqR4bDfihk3dZmeM2EgAtddJmaP2Su
m8dJq2Hdyv5Bu2zeVqrb8Ef5B/E7cBecT894EOtxLAilRSBe82zYeqioFu/VAXFV
QDKSgADSXtgj9c5rv09xQnCdi51VpBWfiN7bBbMQ/26zoWR7juNXB6B+ZA9xTpAp
u/we4wYASG7di0j9ENDwBQkV+TKJzSBU1MrVaF9zm+weraY1Y6IzVyX+34URx42U
klF8hX+yc7KTo54BzIOLWqwAJXuAVk4sD7GohyLNVQY+vFKysir1dvmndwb8Pfux
kCKF5S1Vs08eEUOJDELclL+C0CqE4v9mxoBzd5ZnTaDc+jTQOHyOTwYeJiPs2M39
oFFrRQa9S1vlsjS6DjxSvNRIJdQ9ag9WgQFaUGOwoIQaC6aiv0Zwb2MxeXgWaUcg
4RgMtkxtJmY6ombHF4vBL/UdbPgvFmHhzY9SxeYFqFB8pdnsQCxT07I1zn2VTJbt
7s/9EFzTxwWPQzRO40yNhiq3t98ZeGZCZdvG+qlBRLoiarx9ANvIomc4dYVXzCKy
30eQrKh0yQLkgYgFnHQ5C9Gf3fFrasOuZ7nEA6lIcuPX9HLVJ6zhgyYzja8SH8ja
fONqOp756rqeL/4YxrFjCZimiLhwuwVzYhy7sz2ElSk8RUus9as8aZtUM99dU0DD
RYJm/LPQZpDhY5uGh/QnaadTjFgezUbDq4heK9Wr5x2KnRnwfRguf7ACUX+E/aEr
hrV79oRaElikSeOaHyOMiYAJMTRW9P3klNgZ4mBtX9MGItIFDl2IguwMsKdSMr+k
t9bxxJDZcdZLVRwFvPD/cXTkSOych824/O5zL++N164YRQ4fX2lq//r2FyDQTUap
RcbyhiQZ2+pMXeN9gmoPgPh+E1MS3400FhmOX5bWjiCJTzmi38jeYWFkwvFz9yHv
zElgE4l8Z0vXAElF9xAEMWMaweAywcsPxYSFxDhREQfp/gMC5ZLG36oAm4BD+mTa
szLNOo3GBeXUFpY/UkcONluidTy+yQO9MpCKeghLchYd5u71cmVpzCes7CeWcaMf
l3fvZ2TvgJ0smXZmg/AEAVM8N2BhrikNm3Hd8o2bFxV90w4oYIQf0kpZAVeG2A4c
rMSbaiHZvhJlyPMmDMoZpLgmRpXLSycvd7lfimoylxaR1JlLNJcPUxVvfedRdUJc
sKlu9GPt8bQr+P9PFcka3wy8GzY6Wj85FZ+lR8hZ2GeZEFGDw78GF61glWK+LDnV
ILgrqxlf1KpIoc0fO6MHlsYq9a8k7rf4f1eeT+XOXUB9GdtNczHa7krXmVvoibkV
BtwrYAww+ERrCXdE++4uAh48v7/yTPX9kT11uinn64dI43gRCeE4YMBCMKzcXWJk
p9JRfv4KyUyTAuLYwbIYsDW2L9pkJuvqH6OYh+FGLEFJnDf4AKi5QLdYFUCzjwQd
DAeKkNOupA4aHNDphcIv/aNjbcewWWbUvaUl4J+xRbhoYIbA3vKu3doNJNmUtZ5C
`pragma protect end_protected
