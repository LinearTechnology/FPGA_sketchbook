// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ee4axti+loKQJRnYX/kA6KcisClJ0B26a9fuYIig2FGyEbXGQXYLuepFBGHFdSMU
qanwNgYN5iFQWF/9n2nhIWHtybofJ0BmhqB61aoa1uazBXMWSPOuzLr/1Q1WeGoP
W6DfEkH3asYDt/riVWRH5/tMCM9yQH8AoX0CJO3Th44=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3120)
o1r9ZGSE7ljlJ2D1MxaiFILFxUwDKybwjFNskbdLzaC0Z8i4KyLhfSiNMnN1tDba
bks5a7K81HXm8V4FH8SgVGbIwgeBK2IQo1IDRZQIf5LLrZbIGTRKcnPjUJjg5CVc
EdK/iAPp3SOD3GwLZa0mC+7CbUbr4j2W3TimmBJ5ZdZ7eDgxLRS38/9RM7vaIXyD
eOu2OAsLi5yVIVYndCCkhnSx9j+HGs/C7SeqSPmWS70E238i0YEU9upKMmDk7ZtV
nxe8X2jJbbzkaP93jA7ZByAWu+sNO3mqzaAK6c+OsEILkp2xJB7PD8GLXZDXApgE
CVWs5oN4oYTQBwqFyQxdb0TVbfIPTbsKoq9GLkMvpX1MpuHE6b5K4ddERx/xEVom
RdwsOZSDCjRDtfZKGVupcr1gBdd5LDqVxJ1hWxGDX4ci5cOVDZf97pOJ0XLIujPp
WtOu+nTxJVrXzhLX6PU8VHZyYET2l2TYJyrUHjBzWixDzRUStgCTF7DgVg7obDYJ
78UidGrLIa2JsnjHugw8JALAoS6K9zdajVvGck4xSLokSCOCNNO6+K9tSko6uTDf
5LzBqjzfWlPUU9uviRmTw7C5i07x7Cxznt9l3ala+jnNw1zYGaV0MPITFUsx9enm
7TEm3frdONnktbudMHLM7XASeUv25ib513T07Fg6cn6rvTG+bJTG1x7o1j1SlvnP
aif7NHl+/NqQAoyG/IkBfsYhEUhzlxm940sc+LrrvPd5l2yny6ikg0KzGccDE/FG
cbeqPD8QtEtRxRMoekT2wfhK13zk7g8QqJpvQg+5leSi6mO7nR3w6x9ZxABrs7uB
qc5XYBiLlroqw7j36BeClxGeaKkNL4dbyqY96VbUptP6Xpn8WJvmyf81AKRXyfT5
G7k67AF2b2IVLRgoAnHZEOLe23DHw2wPCh212bOe6/BDxG1vZ/q6YNWWavbY7PF8
Q8gDwX2/c9h28tIxKS8DsqUFhU6T8gz8ovBOe98LD0wRwV1jw9ymZp2lwv8mACWl
AFPVIXm/GS2kjCPDaB7IFWpblVl1/7dhizi+8cwgccDwUYJjMP9LlxroZ9/m/3HO
V9mDXyRf5O6M39Wet04rfu2BpyqQni2kQ+6q/9x960SYJLl6z6y4HuhXHTkxpeG9
YnxSTF1rGZmdzVKbd80QGh2QOnu2w1oDF2is57gULfvds5yS6TQFT8A7V1Gh1RRc
rUAJoe2mfwppJLLLDL4FlUK780bwFDN5KMP7IMQUpu2PQVeb+Vz2uAxJAZf83zPJ
hOlc2cPRhEqiGhz15garbDqZZzJszrAHNfbXz+TdIEkC5y6m0mz/hrFnT7PXSOkd
PbcEzyn8twYppCXc/SjN0OK7oTj60Iq8usfqG1jfr158r0vRgJoyZiBta0Wj75wU
77EsRcrPwlMppfCafYVMpeCPScjB7cgqBwleOID39eDsSWRakWlT81GWkJ+tp1eZ
uYJfa+wjo/jBG9MytsQREEcMYyVW03lv3uYmequk/3jU87OVMk/6cSMDp2fUIGud
JNd87K+3JagheDWTtx0SgFY/3tUc1yVj2ZKLkVRbeQpJSodNouwz8CZSQ/QW8Oqx
YwxqPxjYQ/EvE+CB2JJnR/YDileQ7Tt/SnoALJ7FKTc/oJkE5rdpKba6vn3ZVapp
/ZPt3/aAv3bnhT6VmxjgHmhb9sxAv5EHRbPa0kInAC6Yt0Tt23fkS7Tm1rcjgWvK
LE9g6/9YG8B8rchKT2s4FwzDc16I2+RIXpdfRi36HPhSBZ9CZbveMtj2Fff7OztX
XeSmuicVvdGNPoj4NL5xPLNqwzSoibABx5VEdCG0aSQzb/5Jlx3vXPeLW/9JOxah
oLAScqQHC+2jFYRjSwIp51AUodEQg4wLhlhOPPZ+2t+qZf6Kd0nMPMyQhjf7jBbN
FVrXvW9RzSbsEzT7128BXlZhGNHYv2b6lQy6OZNwf2Gts+TdmpcWUtIETLOkZBpr
WZxlXxW29FCIIkjsmlxFHqxSgbnvAOUC9bJkUQjZ5q9HE+k8XOAYtaa1XNhQeUSd
Zk3eRuhGmjjjtWRY7h1XL3lCzYR7nDMSMNolXtXufGV9DyGkQHW7Xh7wYCuM7wAa
xYDaAcrvJ+xncZsQKD2AkNQ9yHWiqJmlDDHRklLr42dYXyQP1L0+M6YZ1buNf4Z5
ouWbZPA/HvmSeHELzpRmEx2sJpA6AkxZnSl+FSGR82h4f8Rw8tPG4Ra7FOpTUmCT
YfFgpWbtK9RldsctxCWs7l6omKiFrrqbO0IV6Xncmy2VsCjzpjvpV8lmq9OFrQWk
LME5oG4JThRSMrPs6vL9A8qTfEl2CHonc8k0lrmL4FF/ZtC/BfiGi6qNUSmCab8M
79jp2gtmi14R/sP0/7GzHDJqNnqlYNnX2OAkXBYmH7DMGn1dm1b7oAdzSUgfDqtI
lmXymPdvQ8DKaDTu+c5zj/9+c5uWeHqpdSNdISNP1dbCASHna80TQvy6GTVOdQXi
u/6eAC5H3lehNL9NCpGKbJD7p2zvzckcgWKs5B+0m581rTHH2AStLOLGvsSM2i/i
L+2vCMrZpGzppnXBWNoiE6nvm+ryDnIHNDSATlwFC4OvKK2DQgXgsO8jBI+cLst2
CIPiW9O2ZTJvvCkkgQjlMYJtYb8tGZuVAtHeJu4zB9LPEPLPjiAdGdkD6VWgEMsN
SBGUsTn5wp2AQjEreQuxOoXIIHhhzo0Y8r7KyrrfuoMrK2vfTb2FlReoH8q5tuJD
x1iX8B/hZ4Sxls3p0Q7P10i6KwKq6jIv2W3rED7dvUQwbZWkYT9pfUs8+gq4b0YC
N8Pi5O7jnmP/+yJkgLP+4k+VAiinmR1D6cr7NWD6ZnI8vF8NJVffMzyogvmUoi2v
08CK8mXOptHrxTpJhfbFth90e2ZmVoaSn/cF5uLcRWiMNirAaQEb9/CMv5gQ+6C+
jYCl+NWHydCmKEH4yUwhcIm7QfehPVuXf6crbRuqBjMz2O+FUnBuO/48eKcWj4qf
nRrVNOjqkfPbr+y2+Jda47KVR/+P4YfkIpqZPDHfdXJ781fuEpmt5L3oJUQFUS8R
IYosFMMKQg77Um3zyYaw+WSy0+T9c8ouNGR7cRU2AVCawKAK90DG+YaL0XJi5Frb
xOYthWopHa07KMAqr/RjLPKPKK3DdR/2yUoBrdChKI5EItGrmJDdikPmqpMJYX9X
qeHRrtLGdrm4MIAiEp0NWuTj7Arf+HYmhkgCp1aAKi5CYR+Qtuh2W81OB9ernJW/
UR0qWM+lB2zxiynXC7evIYQpzVpCFlsUmIi3H6289DbKIX13hSdnNyScWwhN0kRw
3EDIK4cQ2C+GxxzngFgoxdd0q+FaU8TdZHuNt4jcDqB/Ng+TYZpAJvBJwozjnC2z
5AyZBl9kdbmMe/IA3Alak8GP5S7sTOY+NZhG1DEzZOiLYW0wga2PHRO1POvI44Kx
N1SQBh7pj95Zmo7KTnqFmFWaa28tgN6VMUFZN3ZskSFDMNUYRiQjAU/oj4JlE0hI
pPB7Fjbq2fu0s9tJVvlxb7w6GVgwp3Qy4vY8mae/+BBGC23VlojwxioJcjfzIjx8
usnlGhAyQ9MQSioY1UM9Q4aDmZyrDwCQfQnjikgDdP+aTobskpKLYa3WLM7sN6Gx
mZSdQBA9hlA+0ELFkREk0iR+WS9n/Xhuf+VgFeRIJVCb9BZNMHOuLrU5IonXKUPL
XLXVwJ3naNIGBRjmJT3me+9xRFPuwM+GANgbMfXogjMUR+f2BrVrJ51RGspO4G/H
SoFrw/0q5mWfs39DT4usbLHDMTFe/vKnlBTk5xYjY/A9MvX049pUWpWnKlghVZAm
xW7+sCYlqPwqOhKhYkLLkZ2VrC39Qww0lZzhL1l5zQstncOjOojrV5oxgydShZHQ
GvoOu9OKvoQaQSwXtx7gMpuE2nxoHlD6BhEClybdzzdD+nfsT27OfUxJW3BOZEXS
URz1LahAPXVYzOaqig8s0tbn41R4O5KnxhnBoyjWb7z4xj6mqjLZg8sEK22JfFt9
4uhXdX9Rbrs5IF63Xsbh0fmqR4MVngr+ahE2Q5jVYnxlz/QBkurd62hXkdYNyx1i
8cwDS5HeDIJlS08+UisH0uqORO0xgKLmn17k1izp3s5z6nXzgV16wG6y/odRMIwi
`pragma protect end_protected
