// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nRu+Wrmkr9aSO80iyacTya9anuLaQ7Fg1r65Pa3tlI+c/S+rqPyxjBcN2rAVZcER
5gySEYeKUAM0nf43dzdbrzn1H23aCi0VKLKfyA6yCR6TU3dgbTT6yIwoH/NQUawB
mj7snE+L5A0ohQfi+Ab1lBvyBsgiTO+9hSiYMynyaE0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34608)
jharH2DWARdlcjg3VBzAfDzK8v4gmGrATzPlBKOXJgMHYYzdAqhJzQ9rjOy8XH64
dnpBrH62iwQU3vC4iEwJXvPMPh/ro4caoahDpWqeVzVuBIx3HEf4iMPukX+9QY6Z
cNfoZpAiK+NY9J2GtsKN5mWE8Daitd0kI/5r9RrSE2uAJTstIYEuEFy38//MygRf
vf4OW4k8L+Qh5YmpheTSKlCB4SlZqTW1kRcQ1z35OAQ+IZ5Hpb5NSrg5JgT15J5/
KENFpuJn2Wknu0T2R4M+V8NmnKopljXVCsY1cyvgb4MqVTOTGWcpSpTGWlwVl5Dg
FjJzbwFSH6muB1SpHTkGI0pPK+OyYLoQTw14SVUrn+3iWRYuiskFM2vfVh9pBrse
x5IBYzVUHALY5oVx7BgotPewqE0rjk49x8l6l5WHkm7n7UENgbgQdt9P/sBMuAyI
3hYwK93K0E4wDEiGUySNt2M8wCASEPSMDM5Sg70s3kzjkBXy2XrNt+c/BnCa/CAZ
s61KmdfUa8CTGdNGH+oRKoaJXlc37j1JsHhM3AHVQ+6h+yokAch71ptxyf1rFstW
DcNwjIUWJtaYVEicJnsYWdFf2J3uj9WI0PEWFS2Gh3iV5yxGhpJY22cFP7rrYa0Q
AWFe9qRBaCXuD4o6QQLXgFfR00i04IQfUuwZyVQuyp1LZHc2N1FZe1GZLzSnOG6W
SQ1uVKnpqHHg8V9nAw918escob244GVd09a2dMS7N6Bbcq2XDz30coKr2cH6CaNJ
zuZNYg0/LYoF2jdceY+GQsTwAQxoQul4vss5rgPRVLdF5owCv+5Kr9QiRU0lEdcL
Op0ia18TQa5WWQ7f/+jlK4P7brATUyZ0goEsFykroAZcS5S6ksQEN6HGUTWaGTNz
zn0FNTc/SIWX7/4ktyTAZE/eKu8SD7OIcP2oXfhwjdK5V5hPps6M5XVlIbCYKx+i
E7r9N18GyM5O4n4//Iz8Wrk5sd/MJqOWMSRFcAsPSLDsym6uyOLoWk/X6Ywf7+Ts
JuE0WquOf/VICWxFr4fduVsg1UaumOVlm9P6LnlpmE6s+mGhDuo39+vQUagSRGIr
31BedM0Q4GkImc8jXSEY0qu51g3xLlRJmZWTP6Gjdjyt8Ou5rC/AashMcidVvPGE
5vst9F63luXZZT/sm9qe/XxaEF+/C+jFJ5uikwE5VtexebNpCNVjKzxosc0yPr55
Wski+0aEst3SbXFmmWkMQdS4ULEywCnuH1FZzo7u7DsU0Lwxwlad8fl8+GcXrSYd
+Mhix67vBrW3kHM7h28C5ifwTVrToP51LIvKKMHD65way87QK/Ffa+jCVE30Jg0E
A1KFTgfNKNHeLcTOQ4MAZB56Q28SaDM8jGka8z+gFsZUHMcctYrqkNgNB21pU77t
zO64Xz+sX6Ki0DDzEuXgO6vWltkmAkWRhne9S+K3mK/Ev4JAe/O6ELakNA1kKt4e
Q8mr3gZDRniMyGt/pbfuaZJZhKER7d123/DMH9i2uCHZr4LOequhri+cRkywAPRD
yV0jX8w/qGyckvI4NNGBfPDRza4wtBTBPanx+DF8ChDO2ecC+3epmT9lP0aBG8zA
nnoui9pug30+88K6xD+suU1MmroiHmBuvI6/BMFVOTXOwPbvrlnOWINc8yHxsC/h
vV3Pmxjxy9SOit9GRDk1W3Ie/LZXWXFM4tgbBHaqtdremjFTguUudlTHIpXbFULn
g7eY+M0I7ZjKUzBJInHMgh0RDTEwtfCXl0QhbFM6Xosvddp65zRz967wOlHiyMqV
5wpnZTAIfuLTnvyqCf6hWVPPvS3Z25AY/vm+553FRoO+/rvbwNtnO66AAAzHxKzO
Q0IXlLMjMk2JnEkEoU2KoEJIPS3F73TpqLB+1meyTDkOtulepNKQFCXX8o/KnLP5
I+xZMXJAiAOGBYas64zyLrKIzc9CDDfsWhyU90woASiULYeFLUO0qFJ40abSExOl
00koqVgWFPzLZn5RsTgtMqtuOOT/sm2cTeKg6pjrZByqD1oEguJCFQIle395l9G/
1WNmovHK9HJa3PygdB90paJ8Sxis4rh+oMkPb7boQan8ufFx6/1P5dceSKlors1Z
ZzlaelblBxI+2hh/Ewue/OetoIwox0TAQsy7hyXAkfKjz7yINgABRzUmlK/l2jzk
yzTzGEEm5QGM975MdVU9hXEyDq6P3czmIfd8D4lBf2QP5G6ylzFzkfmbA69rY4Uo
NO2k7SkMhs+2vqnnbXB/sBYA8RXKqp19ygEWWYg2dVgOjIfA1Czlk8mlFj1vKHwb
uh5Z0H+YtDGPvHNCzgooz1Yp+qsEKiaIae8SsegTVZBV+eP6bhjsL04T7VebZnzI
lH2dGRTLWcnUVG1Nv4xa9LC7/DUne0admQKL58geL8bbHOdS/SjO+kLmVB9EwrAW
pUA69PlsuwjCRk0RFPVK0/Ktxvn8pccGhHA+VYOuMv5MX2SYfMhVbytTqWkBR+Gp
yBxsqrdApA1U9BcTOUrxQoQPYyMnrUxZd2fKinbDE29lHck0JbszFt8LeDFu5Bc4
ddyu110hFRozNLKcJyM10U2UZeItp4yitTGYiDnzQNrvRO4se3Pg3vOH/Ijc6je3
/gPngLtrIW9QoZu1yj7cqhtC8ia58zOtCY6+AfNSiMoUoHpgeS9lvCQ3zBhH/Z52
T8dCtV+5I4KMJJPV1BVQv0RIOXA2/7Ho5fgEZsAVM0nM2mQNssyZMcN9cd0sEfdj
Ob+K72fWVF7dNSvwJs35FKeIzEXt/bxZUD0VFaNUuFFL596BhPjdOWzRI1OPacK+
XYlccUKQKRuwaco2uaScHm5LjKnihx9rQ1Ku7bcjUdDSVl2o+LclR2BSBtN6a1Am
B0/l+bTFc+X2bffIYvVj2KRLiVQJnVPtF9PXABPRP5CfTv/K6v3UMUqIp9RY29Nf
GLhUckR3B+ins7kRl92BG66ijd5jopKwcOrjZP6P1bTDEF/8oik7L1eVPjGYf4+y
dTvoz8RIeKnflT/FYQ5N+Si8DsyDfiXTK8n2/yLyXKM4SjFFpS3zHRZ9tgtvKj/E
/W59yyoGvA15vfjPDyGxEgdE5SmrACMqKYvLc2dBKg9Fek6gKAfzahQQUdf/rF6d
Q3T9uxS0w2MLxwj/mPiklWLL60870Yy4p7VBmHcuRK7gAfHr/iMby4iAI3tT8qSj
RsMUPsMqcIWv6ie5074X3JaxyE5AbmDLOOYaA1M9RkOEOPKloKbXBp+25GzpP7yG
ddYrgIX5iYSgKNvhPfwrH9HR9XuXN55FVXbQ5hpm3aNWMfdEdPobTVROR8YgkR0p
8XMlvDk+V1itFOYHP6GzXFqWwQZ1mPujSBKCBJTisVFjMXxMGA+n1FwwcRyVLt8k
lMKRgLm7hvyx9QCUO0LD4vp/NPCnVkYPJX2XdR3M1S9Mz9eMcx0TkYnPtckD4wSV
1hqWzKvVGZU28q0GLfNPtxg0bL0j2h0ptzuCTuFiLdaygSWQREQz9GVCawcLiyB4
e20roGfqNrroM2lWrJ7wtz6xhBHPJrJWQlwx3A2iPIi/+GracUj8q2ruD1N3WeEH
ARGEbfc72gIXXqUaBiSE572DmGbGhBiNeerjNn/taVeB7Ankz0wseZIaoupIh6rY
gy2ml2ExmW2OZL7g1Z1owEKK+fNNIYJHD2DU6oEPdYByvC/TK+lnG/V4Mlsqc6Lx
2HSXNmUJtAqGt4C+TqGRHB1igmzjPtPuI85XVcUPFHm2VjEpCFNZcxBI2iNFuGp1
jVpv7fFX6hwaiNkdVB7xWONOu9j9DbNAM5CmzXn/7woT6kPUOcP+LrKWNpbU+f98
OsLz4Btzx+Yucpruc1GzvAkP4lV4UKIg7aWMlCz2PWJmHNAjOGCvvg9rdvvoUhd6
kYV5EoVknJUonG6LfYvK+6YWi2nnS1WnK/ozEDYR+8gv8o2waxJKkx91oTaFRttX
PFfe/U1I1tncyBz7AeJXv4F2QhfZZNG4hapGvvzXTx9VXD75cXK9pGW4XiMYYMSL
DU2OUl22cTWL82PSt3aTUkd7X4WBVY4Dg+R7FnTUM2RGGiVQ+5dzStEEsU1pqAre
JhCxHmDffAMD5Esyel7cx4d4pIsPm10ucGRkVK0Tmne4WPqI6q7tSKEnavNE40l4
SCoJ0NXLDCIVHxeUozXvglib/NCOF7dV73whrMwQZIdIYbD0fZGgp86CeyTQj+u+
duZdVdGqNE4zG1siW48AeVcRX6Rk1N1AwEIDpdo9zSRVdjAyHDEGe3f6G3MaZL4D
gRljqI2E+QbCZgMg2C7H2xAXHOltDYDDRNRscjaVAi4KduY4dDzR5WzLQvwkWu73
P0SI9BtnhlgwqBC1Yr6p8k3iJgpS6MDH/GINOYUJGXm5o1IafUZwjkTDfi7CreU1
h/7tGD2OlIbUSlGszyx+GeVR21jsyj1XFNXBCtIuzWEqGFWOccF8w2D7MiD4JPr8
Jhl+kQ7ZXobJcC0t1nOzpIIlYAa0GXYgKQp/H2wTU8sp4pYzNSbciGVtP9++u+RV
cMYKZyegf4Yt/EYMw4iYYQRpYYxH3faDe2VRKwhPnKO3MNIrV2hRbKWUGxKFbZjk
hSVajA9muDFoeU/5+P4yNppcY9jK0GPspwtD9QCalGt4VulLoMa1pwwmmZuA0NNj
lQgtBeHU1/L1E0h3a2isUdSL3S892fDPDdvMGusvplpR3Sk9KlggE5QKi0LHGr6S
Z+qb+klravuMaIEV2gugaSD5s2cbAQNDjYjQt/J4i0l5GJcSovqrnq4awKXwHxQZ
3ZJJiKdRzh8N0gydVrQj/0IodaqllfuI19daRKOEuNIzbRwaP9FYXUSrw4QQrHip
FbhdtZtZXgmA5FeqErd/68TSOmM0QoynY8vbw9Q/qSb/77r5E4A1eC668DuPZq/2
sCpshYkyC3pecbKxSuNCnh/rmRs3nGI5AF/6cc+yTulkkYCPZtRijjQG+oyjM0ir
0F9VUlany8+QKoNxTXzqvDLsi6fWOQWL/UWlSBM5aq5qjgs92xpei3IRIB99aR4o
1jiycir6dM8Pgnv0etSKy2bv1W4NmRlAQyrPvdYonBVw9OUPxDCFdhePSyNcPBJp
x8akZ8PbembPyAZsbfOvMQ2jAtGtolialGvtdsZS2beqhlZp/qs/MkrGEKxrhY/Y
oEJCu/mJc+U0MCDCldJdy9Aiqysyn33E2F/XdHdWD1LrhQjfHeGGCGFQnvyvhHxw
Wh6UX6jiSXPkT/D4SaaRcexfG7LsTKbSNzM73SKrxSwMb/1SAN1uJC0lulO0IqDj
XVcFCYcAED0G5Rr3f/Sxh9YmEOoEkGy+v2+JibSfusoD9wSenH8G614T4t+wQQKS
To20wOt5RnrDtjbQH/Jo0hZ6pPe63RZZLMJgd/yBPuZ8SLiDjKQ/4NC0JtskLUV6
ZTfyyDa1Z8035+euhBKo+L3A3/OcBcHvop6WRd15Ss9R9yo+xsKviGpNTaAeBWCJ
kxHelN8WDMa911ppBe0fgj0YP7l63itHUUveGLExfsq8mKiNDyVYqCkeT9wI6cEu
5zkhpM9XB7PqwcFQ6BUfIGqmvRJyIKp8+Z0QZJGC10apQUXIusrGIJsTQ1+TIf4e
o2f21fHx4QG1QNB8ZGaplcJ5yzYo1B8fJC3qmfhWcoT7L4W+Xy4Hnxm2v94FVnvR
zyAMPB1GVTc3DXeA2Cl8G5SZfESU02h5L22aaDyQHwIVrLiAk/JfY3xDvNuG6dhe
InkeTWfOks4qMFI68hy3tz9PawimkGHM9yf9KuLDuMarA3DDHCJQotE4NHAJvDCS
+YzTkEpzocF5ZUlQF/CeF39gp4v8/WzewYn/l5pC+6yhqwkRj9QKaHk6RvgKZm+U
ILgWiqCbEalykfdf29aT2033W7xUH/Oqhsy5xoaCIO3Cc8nr/E2lrx+DNyzmyGw9
8ipMzKIs66+0xhTGt3RO0Wk8vy6hmfWopwCIWT74VOra5d/xrcA5ts1T6F0LWe/v
YObn6HSCxhDVA6TnXpKKHlj67n6y74ce8A8i61dLGaaPlQLAS1E33dEQuUtKi+D3
NfbScEzLwADoNj+VTfxA9aHE+caBJObHqz7iaPOJ3Y7lH27VSuxarWxKmFCam4WL
X2nxCmRUNy1uoGM7lxCw1ongSNAuKTD7XMI6swr6Q1+bhkW5OmiUdmuaLwCdznN+
sq0z/jFqlKDP6RVd5OTzVs9Uej/xJQRC5NO9G6FbNmMTBboN2hdEJJ4eLbn1MlC3
RJYMMDIGGGEMy+TjdQFoD2R3FCpuvMRC5z2FhL4bO/o+nWoBdsRp+oH6SQl1IPrD
3o5k5tHEwFEMpZPzBbZ6AL9yDWUjSnaq3Y5CfyzC0h/ouy3lacCrL8HxySL4qZI1
ooFxkiVvFg16C3BPMxHeAaEtGJvkqoO5JQylmI0HXMP5GgITfD7iDuDzcN2nAdnY
VRTqdU7NmrTTBRXHC0YjCCusJ4LsvF+IPSV8aJ6PNeHBhdd9oIWprvvGJrjyEcxf
2EWsl+lH1324w7ETF7OIddio7pSgSA5bUP1kkHBrQ6V8Un/mLSswyFCRKSvXkGCR
TxgRFA/V5Lap0+L4WfUS7NfHAevuVSMl6VXf8UtN0ZB7QpZw/oSxovhyNAnzn8WR
XH6qru7rm8kvF7UzcNQOBnpY1IPuP3F5m2LJGblktGO6pT5pnzEIo7Et3jsn1AXQ
N21hCFScx+6RokCP3Z/F935TWz9UCD8uuhserizVhZGKWV4cOQKer90AcpaqOowX
XPMn1BTGB1/DVdxGmrR+z1Br1RU9SwcLDdbwDhCo6B0v3ECd1SPW02+uJgd0WO7x
BjVQ1fBJWtcp6d+xIBsgpfjUGP1vVyF+ArRgTPl7S0WQ0SpDvPXmTXGprRgtE+xK
6c0iOlYvb9epl1zZpH8n1DrgETeslYc+YgMrPTQmhNxHTvDs53nTz023slO0SAqs
NzOfJFz8COLSqPjuo9ReqUP7b7iLVgoO/GsUQpJBidhNNli3w63EX0PQ1TOfrGQ0
VmF4U5s/shH3ewy9HnRcDJziV0jh57mFzAxlOeX9vrJCpHdkHQZ/xnLK4U6Xzvqq
W2Kit+7O8I6j9TzosXSvvsGYU5m/uo6wWQMBpzTP59U2dAx28Ge90HEl47JUmWqH
ES67goLNQHLxU1KcyHOim0uNmUThkgSyjd7Dh/VF8y5fMRYItqxpxAMdX5s+XZaH
KPaacbCJywT5Z0yu65QOqylJFpTEGVRGQ5G832UDMO5GF+Ru30wM3Gsh+QtINsmm
iYigui5QFsh0sB/veKIWSotSa3ixUHr4JGmPcvcW/2laD2cNu/RzsJnkiAZTngE6
WCE9KIMy03KJvwRxf/WSO0wKoddPHeBUTXhe/w4+9sBXPTPXHrCm75w+hHkPjtX1
63FxDWBTEVyx0l+Zno5g+SGnM6OiM1U/ux5KY5AtazCcMUbs38AXCVAga4PaHk6B
HJE8OJaKxPo1iH3J2/W4LaOTEF0Oj+pbIqVLum7Fw/Nfa5RmX3312ODWfp+Z8RN0
UKhVijd+H9H567n8zpPoHdnNq0W3eYJuqWyK08sxBiORrKzyGr2nLePJqH9lCpBl
hBwc3x/p1OxXmON6ZgH6yP9ZCeKvQicMmBBSteK7FVDivX/2v6ESp/Jni9jNwT51
M4Fv3pcHLIQUqNsGKjl/FWwzhcppc+gJejOIpOHDL7M/8RmfqFbD6rB13XtyLCwO
dTG/jVpkQDa90bxRIArAaaANJYgPxu5UjT+lPg5U1Yjir5jEzQ9oQo/Eh3WnXVrA
kpj4j5b2nwMnfrfGSiy7vzKnGYh4sr3Vt+nEBqoHsSFr5M8GDL/fLLwA47MGVOSw
iaElHZykW0Zwv6XBczH2FTUZ/YZkW6jSisR6ibLEq/HaEpNhrw6Zg9yN/GJCgYQ/
3Osn9cgKCLxh+GeC8vdJkjimMokm0mL39UAOTiHrpvxe/66NN5Q/heO1gISc1Sr3
iuvNUfcWGXa9aMankAxvV2sZrb0lXghfBhEcyU2+kQ/StCQw4ga0d71tL4FLSbzd
EpZN+B07wSo1KsJFWY4YGO3AjSH2prMG19sq2DPfQ/gyIeDuHy4/mzg8Qu8pj0Rx
BcfpGJGBX65u8AZlpkLaOO/GPMQ3Q+bTfyK4HGoYJJlbbN5d60wzlq4xSbFh7JQI
V9aj7W8RMLczrnQiCkHSITiJHc59vsGdst/8zl8yzqRmSty3l01QsFQu+e1ZyTaN
+jqpUgvSRj7xIEnT4bKhSr1yN5WUHFARfBs9PhI2YuZKvLpxm1PSnGjJRDDXEmh6
3QKvvnjLanWwzTkegOv9zFEJC5fE7+KuV/yj6TdSLdioGEYASpgxh/jr2nsjNXom
PMr0BQcn22omndgMPuDkvKZAYVEk9Edw8BrgOH9O1UKEUWJ5+f4gQOj7LnncXQkv
CNSvvK24LTL2IsyZfsZIa3vT5kdGMS8DOcnnpMg8D5Wdmkw0dmCVjz1vCFb89HaB
8P5dX0TBbuDHdFr+bOHu4ufos0khieNDFKJ8zbapdS7VYKvQoNFnpIfN2UV0SHvf
g0s3+CYXEszzyNQqk2j635qrDY9dBpPJ7bJiAx7NfpVIybW7vDRslBteUptHexHA
Z7r2iz3izbcj56HGWbzqD59iENVssoYOs2PWLodrD97owqugJ5PQCB/FRT3sIzBD
c3OI0RMljrC9U8tRxNZirl6Xon1huBBwvvJi4j0Rz3LJUeTKatc/B+k7JO66eeGX
u9KlqbMLxkbTlxT9tD1CJC49fC0aiDblTX9m/WnCKphR6cUQtiXqPk5xjsG/yrQQ
eL2vg/lglptaK85Ho6wJHzYfMF9LQmH5CG1JIBd7nYQdXjbMSJri+R0NkPaVq635
EtR2yNZ6TPrA868MNaeNpILWL6zmCf6DpJ4unuSWSMz/xUDF8gluzrXLpLXwHrRr
OmAYx9CNQIK+VtpkJQA9LrIRTbZ9guYOWk+2ZIsIjOQIGXjZivP7P4Ebd2WjT3+H
GESwKcZkj1gvpvq3IBHeA39lkFOJM1MrBjTi3TPBTTU/qlOfiMNTaxQRnmtLB4hs
vPQUsY/FCHADIciflFwcpvld9NiMNfc5or6+hOqRQXmfG/EuVk6aJNvitb+du9sB
UQp+FCEK7Sev9+rWIsHKQ7ZcPouwH3hRtnxtaJGe8Ui85PC7FDK3SCDeoPRZ5vY9
uVaAu6gUp84+rDddU8q02MZZVJ1hLQ7xiJCzZQsLd+AuI/PxmEy1FcbEHpaGamq5
TaRAxWizkXE+2jMwcDWekAfkHHd8j3szmX6bU8NMEpL00/gsC6ncWvwcvKQ48MjI
UrfcMvDdQBLLoO8bb4UCjYcWaih6+/xuuIMUBAdvR8HWCgHOGFr7dIe0pymBYzLL
CbrfVZQ/PL5jTjazHIF8kLAcL60Z7I0sTPIPEWaHq8Q8Zwrl/ohME73HVjtPB5GY
asBqgDssF9C5cD90G2OtHM+gsB0E65injpJU4AXen4e2o3RNHTDpOs/JQTnx6RsC
rZjmD6jbDvhP/Vyb9uNciZHrMXABivpXu7QhYt8xuKHpeeAOR3O7zbxYdQsSfxA5
b81bpqD9eTfSxIV8x8RvYi/DB09Hq57oA6XQQJvRZ3ZcFVcN/6xfr5GdPC3n5yER
gopOr9kU/GlAvSHbsw/NG6X02gtnF1Shgk4MCt5gAWIpoc+DwtoHJKJu1xKBXMYE
9Je1YXkEZu/hOnKNJhNuSVb/a2gswaPbx2W23YdR9+5VnbJMqd5qlxdZgzpOtmLy
sLYECK37Q5vRTLhUO67Imc3G0tW7oOq58IHmEdANZKtWFZItmn3rmu7qONCvYtXF
t2QZ1OY0n0/1Eo+K60vDn39aM1TurmivRtmYhyFl1sH0EsfYyuJaq3diE3rfjlOM
5JThir5a+IozADPJaeiF1+MSmz9CuKCjfGcRPuxJR2GVzCepYwrlwk8+N53KzvGG
seP0gvykJcMHA/vWIXctPHeWFB1vaETNK56eopl+pBxPJwQVzD3XWuTHYGNAx/0r
RqZ50tDAsHv3U0FPN0avuL7cyvoy998Si+Bo85FJ+4IopiSMhazYcQmd66EMUA/7
LE3dvoyNDpQplTD8cxXVLHYRnFWAzJzGu3vS7YLuunrKW6+VES4KzPSsDYPMWP0P
OOH1+7XP9uxPT34wthBiIm4u7vdzPS5Ccg83V8q0v4YFMxQxZ9tiJuw120kr9bGo
xxOmxhNWf2IJoNb1bg86HjcBLOrl6FX/IzOPfj4rc2j+nvPV9/a1s4xz+Pvs/QT+
+28PQUh2hHM5wbCWS/l+orV89NoYVWBim42jyQbO7LGQrMX1r8i0AZLjhupbaTrN
tUk5OE8OtMFe/iI2n4X/lp/rmONbVh71zgi05vXNWqgll3om//IIfVe+r8Zg6UYv
MA7DheDdgIrX8cm3bsrJJJtxEI2UHp5mEyKrZk6p6RLvllsHj+Zd5AFksGRqESqO
U6pT2zubwivIBryKsWBW9/3LTtnDMFWNtmBnAdPqtBo13SfY3nXI0798rt+rTYb2
bz0Y+HIU+ctDGVslDAxoCy3UUBCpQ/BzPiN6Qn0nyE4QAZs/WNRhdGNEieMA20vs
AVplshmqX+/zYF9ntUqDXQ/d9hoq4v7j6F95RPDIfkLemZ7PSsMHjW4I4ZjvDkO5
WPQgImB0TqB5V0aRSGqu2r5DSCIdn6B1KcdzcMd5SrRNLkY63On/uGLeADBmnz14
ECw9xTcGyqiGd3/FL02vH/lXAeD5AM/POueXgxqcaBLuPH8IaRlcv2EP+A15fZk8
aoN/E4NSmK46kktU/5Otzj7kap+2J7YAFZSPZs/gDfKvBL5kyxrI7DmkWkgMqyMq
rhppd/hiv6csUQf3SeXpjc/PTDyHSpt+fQW6HdE86WfhVbbWWYOOUPXRZAK+ik45
54WmmBCsTJuJPV2zuQwbi5qwGCGv80fARJIY/HAqJaZbwk3cz0vsf/DqqVs+TS4z
R71tLAJ0cgk9c7g52YQdp9A1jj3KOArxwhA/mkh+mST14NMFwkjbAw+1zKplaD15
yYYK5zgo93yuswYRI092MM1MuzkNyRiXv9nBqDTGt3w3MuHAoDr9DxO3fy08okGR
AFMTWZTOXiU7qfZvn48D2X97h4b51iz0NOBRI6yoXN6Ow1xAaf1+yvcqEfs5mBXL
DETMpv23qGz4ucBW9cWxMgc2aAXfHFZDa/2uy6LGklcVKSUAhe1jQ000VeBjdQuF
m5iXc5cZQoYC4hl+ImjCp3uzPAbE8X/XOdmQJdb2GLwA2FBWdYiemauatbO7d9vH
fetzSlbA02zwVa6IDxd8cmCFpFEfv5S4bfNd8tatOpfPObZ2xMGPNoeRiFzyY/Ij
Tj/rXk3PaN8nkISUsnWQr4hM4NkwTz2fiHqqbReW0LHIOy7jeYgoZLQfYAOkDf+1
vcdC/XDTUpnFNZ9ltP/Qo4mRWLkGjZo5JJB4VE2AYX5FZvmSv/BdEQ0efGN4hsvt
Poa4+yusCz42elnjcR0j6aQLm9FZCbQiJ7SrKa/erUKvCu4A7fEtnohNS0uHhpIi
9eFpWa8fWJpTPikysWvdv/Sw4dhdCqCv7dHnMMDUlz2N/4E76klRVrqcTcsyWtRx
2QK0CxiEutCKpDD2q8XWoQ6Ag9YAVwELuYajje8WAsIlgOysVVxne0Qf5YRl0VqK
jNSmsmAaV/IYca1c6AcwMcQMi4uC07unbNjvAp30MxYu5+OlTbT34JwBHluIhPwc
S744TeFwqYxffAm8VwMi9cbl95F7YQHEZXXKKsJpY278LgLM4fOmY7EsROjoTXqo
88S1OGKGRkBdpEtWn7OKusomA44Gvkg8MeAgaJfmOU+Ay+U479qwt72Ks9bQcKcM
FE61M8NDmCrQdlSqc1T4EnDyXNGfX1fbWIc/0/EPgU8wqw70CHOJlgVLE4N/8f8A
F6hrOL8WO5HUTJjwqf3/pj9uwhxp8FAWYUz6MjbOAml72rkClTwttvsBobkFgaaO
NtNkPhNasAL+f/pz2LyqAFpk7etT1z9Vqi5NMawkrTKbkt1FKIDP2CZrOjjpsV6/
nmaFjf/Hk73Gyq+A1ICgtxNAp2T4qOhwbQJaZjQkG3aSHycf6aSJbXBvea+N7kyX
QAVZ8AUJjvHpW68SBMDxucTsDh38/s48zmBuLfPL1ZNOBm1DfYu106DNw0aZULcV
/ep1s2VDSKscgrI8gHDs+1AgslquL3ZcTModvl3YDG3mCl9wmTh6O8u2b8XdWCHs
kQJoN9DUyPe7v4E68I3O/6zJ+HD5RACwVyIiIa/nLhqmzkNH1MOPAN7qlUMc0+0w
HbIgw/D1SGj+nda1yUVVCY/foVEYzLurlQ8YTVKKwcfGOOaknIPtDDqZ2y2Uzwe7
f/uNN1f+TMLozPJxe1O5zHW6BES117GkIelNLjAhCDFy0bNdalSem1R2h3OfmNdA
rpahhboNm98STG08GT3ZT+qALwhQWXgCXKAB1o0dNjimi8nR9y0bZj49tygyHF4L
vT7yo6j+md8RS2ytRByUxMjFl5Uy92MRVSgYVJ7/DBMkKboTG3X8UfQNh4DHKn26
G1MMJKzPVpVVMaI1jUkBzB7KLLdvbtAxtHKxpWv4GR2RzGir/4VF+Pghqs4qfih7
UkaepAPQ1l4Lt/rpOevTCCE4bCx9DO3z6jEPcvZ6g0JeE9kG+FvKcTmdDhKImJ3P
CCEpAWvzOUA0C0hoqelQPpWmN0BiQWzIEdM1TT80C9XlqU1nQefcxFJuCV59Ta6w
6ripT75Yq+P/H2LwENuT631+n4w5Y2MBvlryDlkSFmSc8DVZ24sMiAyPG1gAN7IA
y5NdAzoEuc84PuDRIVOp2o95UJgDlV/gqeec9nMbui7os+KG3yy9kna+NLOjr6eW
RDxXiNZCblY4ReMGx2u++75EsJrVnQGuPqW7QTaFZdZsh2RkBPF2bDrBndaj3lFL
vLyYVb+cglVBA6XTuJqOakQSmcTirQgw1fCH94J0PpOo7hZO9Ecz43NX9c21zVgT
bOWozp9eOWqfBuFRmjF+4bGFmT/7BI+6k25qo6NurDz74tRvEpNLUGDdki2bl6La
hCZM1pZcgV52fddl3Nl8Ij9/gcAgkLPPpzD+4U/ZA/RzVQjmt4N/RxLp/9e6SRL/
j6sWtTPRziyUYvvQ73yBGf6KBuM12+usJttbi4Xc8PjKCiENsm1EbhbE7v+BeHsn
81f6vf1fwdLCXjKKHtCxOR+oBQdHt5PnNCx26J3wapvv9yisTKQ3ADUtICoNoB7r
3jXcIsM+5WM8BcG3/Z7kaPyVnzabdEWbQkv+HK8f7Dp7TP+5pl+zfRSUjbnDne0N
itgxKCJQGkeLEl3rA8Gm0JjLhsFFzDw238m/oEqlmKdmUeQdj1YvYOcfUxXwW2O2
NCxREoqF7dedR6iIi11km1Jesih83/TiZFObhWvbfn1aiE8sw5F4YKKO4/RfkAeO
AZjE0tk3NogE+NYwW5nZ2evwHQ1auyZTQYGhPoQH7it03lUDFzsBypBFpTBxGCf8
TylftTHmnjc4TtQvwiCbxRGAhlqnkpKyoWqX0rziltpjKGLEjsGH4j/GtLLnNeF2
ljMdzkIxVrFRVZnQ7QPo+J8Paf2xO/Mjzi+jqbhE/YmiRizh/l3tTYy3y23XtAHQ
bhW/VP49aFfXpkiCX+2T+1arLkUNxBJVIjq+fGIUKEYiKBVX5xIe/l60HgCKd4AZ
Eg8A1DqmIbbBfxeMsf3dtiPx8RcGguj0gfcyJ78oyV3V/v4+m7HVxzqFNk0WwSqK
yckWu3O89plKPmoqEzeEQ6OL0YZX5ZPb0vS4Dh/SXj3lHifs4g54mM6LOLrSA+dU
0g5T8ngaWBKkJybAXy+Sm64V029yRN7xcPa7S/hZd5S69WGeJNTCrER6M76wZ8L4
/L313BXjrBcXEPkz3g857lw6CUKDeowoxuh6aZ+fIeBwy03kPby1CsRV50Q6oUJW
Fn03gRK+twfasE8BlzTfpbAUkBrqHxHV0BxojGCX/mT46Zcv37ZGTbkJi8qsVbTC
XrVUDPXvYasbcCSR4qx/vUelwmXL12gr/Jgg4TL1hmUvMN10X+3i3SvqJFwvVkX5
Rl4ydCwi2XWFbWr/Mzbfa946DW4MK/l2xHPXatCxRPUZe1LWXeI4azfgfNjg7D2c
/wD1tQnImmAv4SPHQ5jFiYGJTx5jAduujz/hHNwH23lCxOjzL1HBd8T3ABRsdw9m
D2sERpDH71BuqcAC1xsuaOL9WRNyVxVZJaQvZB0W0FWul8cH0PpaG9n6Nf2qdxXZ
L4n9scD8EqaE4f4iqeZdlrX2oPOTPgyZ1hgkI15C1Z3RtF9uhXPDhc4vx8CxITss
YY8/z7QJfiG2Srh/ve+EByTYLKjmNTsVgExOMYII74Asvc9mhRUPaFe6UjK2dtRe
6X3F7/wzAjTMOidPn5DmwyjPQM/KEipAZZF40ky4P1VC8geBpQbKX6LNhK4v5vfL
6oRM7DTxh+8Z2x3cLCr41Il8z4Vgmgua8ZrIit9JCI/HdEAa5ivKF6t6OrjOApmb
tGvuBSFtZP0726nRRqYDRbTWRxEZ2J3VdnTRCbPcn74IGIodiTZjDRxckM70vJ/M
UWqB0l8MTsbXSjVGqJP0CvgD6lgkf0lzKC4qQAgrOwKDNLsg4mAwEXEg17LQHcuc
z6LUn5mVgzxDf5/i12wBSvum9q/Pz6WsojnAyRNb1lb4Lh/Ldnk5X2/EW4Lxe5va
78WdwziJnYyWE31mu0jTTVwIMCzLo+2yc0CpSd4Gc+G3v58jPrHD97rsS6QQdrR0
4VHRdpbQS/kXQXpwO19YizyPjpjcN0mtUhhdjvP0PwVjDmE3r2DHUsYfG+JH7xUi
YGypLaXtX7brM32pUcfeUk5nepbXIkwe2itVvJ6jbp0l8Kk/7Qi5Z7G3FcHvXyvA
8uZUxntQkUe0+pxUOPCQb4nD7n6V/MzfnNqRpzKIO2edvv8NZAfn9W0lLDDrGJU0
7Wx0zFWrfXc4zEoux4z+gdCdKxg7yq+mBh+CTb0qakDrtsrW90vAcpYptVMmc8UV
FMC576Aywes+AvtJu/NUzCBe0cy9j1MUctLCgz5KhiKc+I0uUkJUZ1TDZmGgGwzg
qwFkpQWGtnI1v/62VaqeMoiNswoKVEcHROkh6M2d+Pwrn7OTqGXDguGa1019y7ra
GB9eg2rVQACQvRpOtLRbJ1mRiDYwh+ocgQyizz5kLEdaBN2Bvhd+64Hll9tBwlsK
noWE3wCCXYi1xwnjElW742TXDu80WApKF8oCfgcuTgoO2/ipQkFPiSdIAxmSixkW
RHtwjyeRRtVZwbf77vkBYhmUyw+AXbe2/+HuHc4L9NNF0Cp9z3iErSY4WCBTD53V
rANQAQD8bKSMg+wBvaWHU+DH/Ad7QTyFvPrzn7rB5X5XKEwIdM4lVfUrG6/JS4sR
Ic3109+x/fsUI18GoGFRHAR/r5w5cZxCYt/aVA/txfr41nCnpOjQxYCiuhLSVfq4
ZOh2B2VzYjQvmZUfuxJJrPTVp9i4JPKnVPAbJ5mPAJz0Ko+Qcagt6U8wwlzBuMJM
+4NXLXjm3nlWy1e1TVU+1o2s+FSXSzF48w5rJbQcTBRNqjH7saNtl+kAFsNUKijY
H5xoQ3iGMwxjrL6MwCK1fpTNAhREbeRCvtkxAHAJIzO/8Y9nIUNwvXZIb4qSQ9Gt
LVqvM6Omv1KKulSTuSXZGFNgaTZ4u47KgK+8DDGl+PHS1abS0yPqel6yhZbEOJ8B
cCLJ4EsuzNEkbCPGpA6tz6rTfVPm/UQXzqBmQaNXWKr+rL8TqzCpJBEFZ1EnWyjV
O9e6uwd3Zb1r5F2vIvS0nTJ0TDEDjR0T8kFRAZQzygH5HPYRJ9mhKL4ssEsM3BtS
LwBCpz9bwppG6Dq4ZHZhbcmCmmqofmt+cMR/aZVJWF0cVVLOhZwcNWApPnxs6C6o
zWQqiooxuLrGLI0fnzGEH/XjSrfqtWZGodAG6XtlVyi2QQqfxkBIVizS506oUz3I
jg0g2RUlem2l/SgzBYbGK+oifs4pxW5X+AHk9uxHrJNEheUfM6od7soVNg0MSX25
X1ixV/KqYv6Oy8Z21D+xtLvgY9ll6irF2ct45WiU9ZDHIYMDcL6EPNok84+wHam3
VYDaMB1RBTtCnmIAtBiD8Hgrd77b4M7LNGFZ0A+nT0xdEXG9SIOGpTTgp+xZ+uHc
8dlEyY9lVubBKSWlsx73rSEhyHvK4cQcOzi93/Cqbw3LRs2tI1+EqGD+PJhh26hj
H1/kqWuaeKRLdu+DSFqHr5MZNTq5o5Vu8ap1jxAc/YgogRM3O8F0WaL0kjbg8qn8
DzZSPs3jf13AsrpKLX2c5pXngt/Hr0mgTXgydGmLJIJEO5l7FIM1qwjq0gDcTUD3
3nfdtbRyC84vS6sBu3XTcyL6s9AR6alwhaslb6wW13utETPB6ndTlMQjMIO4X11d
mDecj+yxYZ0D3XbtbXM9zDRIXAFLv2hqi8Q3eQvrOao8lEddbDsx2fWjobo2sX+e
rhXTEdnfR+jK58W77K6wgEtcQP5maa1FwTRYxjADXLDEhXDMVZ9X7aNgUO8oPLSE
1M+uGjG5EBj5sycfJlxA3Y7kysOV8Lc/xVJk6icncNu7+sTx2L/4YXbPiR08E6z3
AwZj0VkkdCe5XfdAlHtRvz8l3lWIPMrv/IogVtB9Ic4XagL/BdpsCTHkuvdFhW77
GGWWg8Ewjz34f33rxXNE020eJypPcMGqpgqHQQS9M7fbdHMeEWOq3w/fdZRgU730
85qDM2I30NFxnVqSPJSqNHHYUUqGTLZkvhT6L415LOVjRUwUUHO0lzO4PiWdCrF/
A0XWnAzeEZ9hu3zjJokTF6KRKlEVyyloy+c7w+mhAJ5PRl+fzcfdudoc3BVD9TeJ
Jes7wbQn8NpSujoZmLRbfzzNzi2UrZKXD1+xQlsiU+05x7o/jIxtx4JMhxHnz/VB
mu1C4FXuur3rrEliaGShTm4wwBDBTRX5PF9nBSsojOgcTQHhbdw43zI1xWLFXD7v
Iyn3udL/J9+avtGfnnWeAybIE8q8QUWgM8N0ofJy/jfAOmN3R92N0PXILkwiestF
xvpfqqHSL13W1tC7SN/fVjK1w4XMmPM7PCO0e3BBO6c+9/ZsfBWtph/WXUJFQKdZ
gLLKXgzO7MdWzELIcQhyzHo8zNWMeSDhB0uformN6MRgHZlWBd+FfSV6xgB89T9j
fLfy9UAiKn2bmj4FpaSPS3vJTy+1Yqah6bbdsLY2SDzvqruXjJHmDFZVabzxjxx9
nO+KcBmTuA+tKJDiGqc+4hVctfaXsTYiWagFioQfjKGc1Q1kXtldd3/4aBdyyGYx
qV3T+OPdhywaXYyWvL65q9o6VFDbIqMr5PPn8u0DNWc9SqzbOYG6vDYDMX8wyW7P
fwGmYJrr2hx3FobyTsD50+0M75e9y3wo+FqHp2A8rYa05EZu+Tc2U2VGnu6E/ngI
CthDu8YjQUzXCJhxR+bPFds9zmX+qKcEdRInSSBCX4LvIxaFrtNAcugK2tU1M2TP
eO4Y65eahV/0aT7FJ6VawUFOl+x4lRzuVQhT4ezvjVY1U2gIZDWfbqk83/fbPSOj
NhDkGCD1Ujfj/sXEhUW/IXi5OhoX5FqqC2VM/YTUKwKW8Z4+ek/G2D/lh4uImNmg
nPnpimaMgSf+iOl9Zv9gh8ZnWloIiWv81rjPNvwMVTX1RIOT7nOeONB5qv/V6jUS
C6OvzjVl+k5d6DmnEu0wjSBCPtht+xgMoKeyv2gSATwmPM5VBZlrfMVto+MHs8rh
gKmwM58uRntuZvuAtV0w0E0TqFmzUmZAVBOZKt69DlfP30xOc+q641HhW4AsaPBS
b0NN6mCsiTWEVzi+5Te3KeHxF21b7ZCrdCM4/vPIBzbfTeHr9gG1908471IJAJ3N
sQo36oKcaMMsbLzmsYOuQKROCVpNcVBEm8/h7AJwoigUMRh4mIrVn6gj6t2OWOuc
C+hwTmNLV80HK5oTxofjwT4j3Uu1jmgKR3yLKWK+AvcEo0mHz9A94aojfjMkG0SB
4lhrC7JKXoFhYEasT0qwRv37to2f8BePfL4x1fGcBcXwqC/7Mvn2zl+I3dveC+qL
IQHUGIXvRuvPsJH7yXeWGOBEdpDW3DUJznyTFmzPCIgPcxfXH8Za3u4eE2emdk2y
Xq9DNmrT/f45E8+XUyenqxEGg2NqrUAxg31aliXFkkDXrTp8IrlwDzplRH4u9xWd
Jn5sv0FiFQNEP4TV3QY7Jm34YBy4EyyoaExnF66BKgt3Jjou1QHC8Hbg/YcdvYm7
8mvsXNwDJoj6BlSStk5A0yiTVaMFSNURTWr3kR4n78OO49BoHQVGIlgkmHY1jNH/
bqkB4CqrOt+4VX26kaKBS780k27ywMpDtiyNpvX5E45u6sziGt3W6uUWwMQuPmug
DoA0ACvCB2DJ/Hum3p7T+PxuElIblpLfy5BeL6K52b3IHQ21oHxyjkcIc4ciVDrb
ApqI5oYV5HKSgb/89aTwU7EonPEINWngBs8XmANcsR1gpvPq6U/iS99s+Oxkeoj3
AWow71uAGsYdhpfAibyDkhnXgfX4xUYnxKcqEjsitnEyjib3oW0B9tARktWkozwf
ewxLV3D+pPhTkqbiXiwg4vdFiNVW8dfzRj4YPgI/gWrgtuuWCwAp/8A2ZJbuNoxH
Hnz+GVmCZDKXp8pdlJ2wnjgHfSWokMpTdoL51Tiw78FfAlUH7KgD7JMOIhstmPU9
T2CnVXP2RZt/0uaqd3kzTVALT+Viw2iaJbQHOWkEE+AtHVPHyL5F+1QGIKXOyk9O
XX2yLheQyr4b7hfL437/oE+dajeks+wMUgnTNdBNrggTz19A/zPeztSrAMtvWAx+
qtUVxT/nmPmvp0jORy7VhQR+cuq7aoVAYozBTPPYRbD+3oeTvKkZ8bb2Q/+VMWr9
ZgbBVn0XE2NRgoNtO23+NnpMvZh1fAsND6QG8Jz5AIoeMswl7lWW6E7jxRdU2sBn
SU2CPZdAvsHXDgEXesDfYoDrvbOM8jBq3dQYxtCVa61HuyJ2RMix41tOCXCZzlXn
gzVuS5OeKRmqh6BLmnNS40OT0YdczWuPYTzG6gqx6eXveUF2XcxNs2zg/9GWDzH8
Bl6Hl5gjLck34t1lXj/v1b1nBLj/r/l4tLySgFv+pB+WFGfamCWeQfrL0Cy59112
fbcHrVgnjJhTN9d4uXwBD1GYYppfItAbUfJUqXVoz5FwHOkIxICa+tEEYXo/RSTS
tnzm+3OfA0tgO5NbSLeg58ygOvHDDPLpkg0NO5pL46lnaZCfcXn3dMG5GHDNgQN+
02VhFJus9BHQbdACJTszA/ZSZt7ZTmLPKfeSITjPCPx997qgFrBNG+bo94W7mCkC
mP5WCb/evcdYhgI2AmSYoUFIHD5fY5gs0OwAKf9b+WQ+5W/+DLD5YpGEhH0Ls2Vc
HnlGUGYSeIiCPTAw87IhtjgQiyTQpfBD/D6sT8KizNHjzlF5qU5wcZcvWoncJXiB
jVQR187ITfsvJBbsr2xuRPafvdXYXZD5Oqer3GQchkeJ5hKarWlYuLh/x73xVQAK
4ojUDa4CmJOUfIlRB8gaqlelbgNEBQlu3MKxHjv6sXfzWvArAVKrVNmekRTeRTlo
eyaHhrGJYtDc+ildTzGIxYVjvcDtzJND/+b9j7XPGV9Rd8846oVzo0O8f8EXB1xd
VHRxO1jk7P9qkk1EhlOdxKm4qsASOnGSgQTOKy9yBZWxMbyEZTwi+iN0OWKGiUww
F6zrFS2IFKXZJuKDCwSiXr1XtSmgaunWuuyOIdCuPD1xv5iQUJIhHOBnG/YHJ97x
29+ecbrcXZJNGEGOXTZP2KyBB2LzzrqiLGcKbQ1PVtSxFP7uB84lsCq3qLNfc1lN
RHGfWfbB5RvjvUvExGJND5vSSkWgMmg0Lhv/oXl09eIaEPEkS28lIX3u0HU64aWF
SVVAHF9A0y2ljG/Re07j2iwYsN9WAWAGeukQWt8RyIyMV1OBBLtapY9s6OtmvGcz
5mBJ8qku4dqYjd1hDJkUk1Y12Exs4ffNxZb9WFcNFrDdadFmA/02Ufberh0E1iF+
jhOsnPIj2eDuHLHumCuujyhLnkkSkh4jsGxXID2NiIJvkAtkOdS/eKe/Bnqm/qZ1
V5PdkUNsJUS36xUwVYukobaGUvOTclTo++ZBWtDZaItE+5ekIv1gZPd1km++356k
vLbdRd4E/0dn+tCE1QX8avLy4haAxT1dSyz0ocFqxjYZqhoNiDb6eiwN/KDebZ0e
sCdey4QAnGJyuj13kAlzpqGiDcYwOuogU8NESugO9mOIRN+UYsfj9mJEJ7EJ1Q8m
5efCRvtT4B3/de3uiV2iDlxK2QfRfognsFZFUNcQr4EmsWx1SwKfP9arc6bDMQ4s
8HSe0YbrEt11gRSbyujFWfRYKcixw0IUVEHTt4wrtALEauZIKUUO02XKFlPU7ozs
iQ24rXNAQpedCyUrkmFQhg77xbD5HgeCjAckph80p0JswYAIuQUCdgCUMa8kR0LZ
m4w3xZjSf4jwZFXw2ZZQN759C5fTwn9PYykNnbGrakVa/z2Uosdk3tq9oylU/3GM
lj/hraEijoNhAqMrnVxSjYKdUokWe0LoFKZqTvQhQ7RsrItXBU1YmMYo+qDjt9iM
GQFvwX024kw0KefIU+/tR3r30oba7ubATJgPiGWXSaq0eYxfl+O2lFYaxvjX10+Q
doQkxoM17g5Row88yWC+AsLuH/ZVjBN34Wbqlvq5oe2ZhuSPNaanNDmJUC4FAaEi
ODYyO8NkRC3rrk0+8UllAPRaU4ocDbkVjfjwVKnSoYlj8+ENeaitdvAwpwH90740
TWyMfCGt9oMdjrWrJBFFAK/cOzPkX3j5NcrAAbthBnVdO3dOKr9RTmfdc2DpWPjt
lJh44hs6RXnjC4GLoDOMxTMZ+ccLwC6B8xaZsocVUu5Px2Wb+uj2bgvVbHJ4Z7DJ
z/rLUbJbraVU4/1uXJ+yJV0Q/s8B/YC4lCpZBR+r6QkWyZnOTTe8IPDqM2NT9Ee+
cmdFXd58vjwc2Mqjp+B+Gat49i7A6qKdQH3F8CLy7rxu7n1PdKqlQgFf0RYCfWm/
SPD2yV01x+70v7pGUpSVHGXgd0PUKsZjOXX1WqSTAjwgdvOFO61mtYsnR+kcFjcM
lswn6NgbKKWIqnN94/4SJeHzAjPHs+M7CGtxO2F4SFUnPaHrxBb4Vuie87CBcdT+
z7N6mh6/OyYtZcKUDCeF0LOvf6Snybm+wNAg3aCerVBnisqdwJFxNvAXp3Y5HUk4
jo/Hl8UXKzd4l/Z5S9EczKoxPAKcRo5mtmEnJOJDRft8r8PKxS4KLFHFxc20um68
HFVyyoGlq7fQFFEqFsCCWXkvkUYErrOXhAhJSY9nKUDjpWUY4WqHEfGbHUbVdPtA
TXq2NLs0q9a1TlcvTPZ7i4XewNY9+u6RSRVQL7K9L5w6dndB/OugSTzqv15EG7YJ
waLYnhWv78pKIJenW579F695lsrOBq6FGuaWvqYsTmvWV73KDTT2nBjw8SKt1IdQ
MR0zgXzNuV3VwUpAPnAG6P4v+QjcvTWxWwgz6mZ0bhoE2597nna/ngEGBQKb6udG
JejR+vakuOpfvBpYyTsGLajiBOIVz6Y2mEHORYxS5Xeb6mgOaVDJaOunoficcmfL
MoMgCjs/DOIqi5ZMHKIcB35EBMUChtiRMJHq8pBCKjPP36l6ZAUzNwx6Yw+ZW9ba
rSHQsJi252dMFeEUy1gRcUNq+aL7yr1xfEJoFEhC97yVFz/oXWWyClIx6Oa+qcum
OZZx6uTMRjlaWPYaDIiVmtvIBNfToMjScKw1XZbRIBRA64gKbTobp9gRdMRJFaP8
SSOUUbpae1r5D9d6SMS2lejhfF8WMWDd4K2URrrCKmX63u60e9cXGLwed29/BUVa
muv6VvZxj5TG1HFajVYgx44ZDbrlgSFzlcvvwO0sNQN430IhlBZTQ+Mk129Oq7Pv
Xrkf2FynYQCTqI5Cdo4AvfYNmP0P4Y6XQWg5R6dSkFl2j8ITCYTesL4o4Dp0hJUJ
hdIuGmftUv+rWnYU2x35MXUKnAyLYYX7F0yCDYqzJEoO4L6COUNM4/kk9JL0hUop
R6cMHc90R67qYYMH7RRmpxxr/iPsGttTYexEWkFQjGaagRrJpck7sLA34iN1jeob
ZQDLZSVX/EbNClWes6aCGAjbfuJsHpDZWowXH/RkVLp7IrI1YTh9WItpsWDfXkEx
ytajBd9dpP88U50hgJQ9uL20l0he6+AdH/a+tTpGHjkjQeOxJ2XKAc8EtmZpQjRj
Xy5pAk828c0Jig7WBAe2AKlwyyHSAvTrCxrfg8Igd1YnyBohXYlDNoKQXVQttYkr
hTDldXAffLCAh3p8FCMyD6jhKppPhI1LZa7fCfCc5NOWp9hXi9qKKIBi8idWcGuY
McHvGiySlGMvWujfxl11gYiqqG0kYO+Ty8RPa4wL6hoN+MPnCWUK2ewJa++S/40c
FmMxg69ppkVa57/Lx1fuUXAsW3vSajtO18l8wKar6lpchPA7ol8yHLo+fLVWOIdA
T273Ho3F5iUiwzi9kAhAc8aoIDo0G5wLcqn+az0loeHcx/UlskLpz9EzjeR6ls6/
pVWVk2LMnoRS1jJw4QY1cTdi9ABZA0B2siSK18e4p4ypBabcLmKYWW5YgHOuuAX5
09T/s7v/ryHjp9sDq+DJ7aLg2BDF/Tei4eYY66qgorpXnCk6c7jCATD4J0hxjNSp
V5K7ct5VXFGJEWqoMp4o+N8i3Tye9AuNsViP/7nXvHDRDQe3QOe31G8BqS+6w+UN
MN/AFvsbkYo3hwnmvjZuiSImZ/uSwKmfCZcoaXXe61Ej3iu/biLs463bdLuTHAIC
M7/ssGKV7DFvAunD0RSxy6DoTGA3CxJwuy8pplNxkBTozKFPCu2tjGl7oDPEbIPT
5ao3/dVoRCSSiWSwaYRIPPlepe02V1bPG7Izk1Arnloh0Lae3sl8KAJq+GScu4XX
G1L5MaYLV/t9Qld5Ny7IjQ14RJYZwdY7ZtmxhrQI9myZtWAiBFfNyx6yLym1o2FS
e4q0lEYaTEvM6Qt0iY6xOWl5J0jFGatTyFIWXzmfCebnn0dSxbBR4lVxGou8Xm3y
umTs6EkFnn5DV2tCM1jS/NSFby1J2ubeJ74pJIjueWpmxFd90NkO5kfQcdIaMJhI
XC+lXEzeALBHGyNJu1QcyMJcD5NJbD6tDSsLCDEBGTuT1T38eHCJTR2nlLqf88Bp
M6Ih/adNdFeg/iCsY0r81cfmXKKbPxGZ9eaH5qu/F8A8+hJ3gpbz9bbXyMrLJaCz
2R4fp5WTsueQvxEbHx3l5tmdtqkW/nLdUrvmJhbUfJ0wJ4DoCRBeaBL4I8xO66Kz
k2m0rMGdAfkhhnKaNjgdRHfo8dUE5j44DGr37T8fySw306XkVFFo31p8UI0tuCGz
yht80LBGLLWYMIVBm2STDCOmE2atbL7zkeXNcUPEEwzkrVU6o2QTTOCnoVxPgroN
i3gog3FrqQ/jXrMLGT5al5CwnS9JsE2NNr0Ny1SgxY/meDxqDbFF+9XzeUHf8HXW
LI/EE2F5reh94WFLKHq8Ybz2yPDtZRTuCgiaRszZ7rG4JYTceRqGLPTw67q4mkzO
HASHNVUadPYmo/G97PWqWshwfCgrYurv3raGW3TfuMYUyaNsjA9XWldJczTH0r+3
SGZ3aHshM8CvMXCLbcBEigB3sV43XyCBiLBIJBjz5I/vPAn+8pou0mp0GbvA1ZeJ
z5E3fg8+IuiycTZ/6BseCPsuCdW7HVZagMpLWIWno1E9oRWBWpjI35YeW2Wb3l7D
R6F4PGA9/OX95fiZOW6wijDT0KO5yIF37Z5wS1TwGL8UnmcyA5qnocAzFGPES8D3
ZOmD+mulF+4+AZSwwDc6sp1GK3JVm6R9HNZ5IrhSGU+Mc8ZxXS3BPmtIcf5ebb5W
DUmNiEnrzhqA7qw08vQ57bBta0f1iOkbsVVt3lER9hKpt0Nrsf0x6sDuOf1/jJYZ
wZCLugEEVdEHsmasIDWz9SXosp/mFKbJvZ73dZ9TY6zaRa7y0tJveke4X+xXEkDL
a+KAUZPWV+XOm3ESucUfjCkNQ48o4U8LwPuPSE9XuNkbjbZKZdBeRKJqGow/xBK9
lKxea/LGdHXnW729SdPDuIV9jicRwn6ltQPjBEXBc9v6JSXwHgH9j0zxv9m36zxy
NQgc8HuU2z9azhJgOgE+1SqR41m23SW6SonHcm4i+sd1B02hUrQyREH+2kLkrwZJ
Uxq59RRaidp8IYSlOQ7ionU16UYls1TsAORtDxUuZto0npwyIZyu3l9mAPpEfE1Y
7d6KLaot77BNwLSmuaQWpY2zH6aNxMBN5aRAE5mQ9JfkMmksGmrxtTlHGHqVWOP4
88HEZbUQ4NicRWQ8NWckaK53KkqtEVVmYjlmD7g8WhIehvAh7LPS/ksinNozPNau
BeQago2W1hf7n6tm0C2W7aaoBf/hhrtB3OcBmzpvkXOlk7230/JNfpv6RM6dUhbj
zLCQ88nhwb/BX5McHl9MkN/O3NiCQA3xzvbhnCGuepbWZmQhHgZWfvqXyOyI/SWh
NaVg0ngRqojl+mtNMlAKBSZq3ndY11FktHRKMKYENwAeJmMA0R/NuXcLbznTkHG3
bk1MRvvUJJ0yuwN9ohrb230PTAOMcULo0MHU49ZSodtxoAFR08/85FlbJjNS5xLR
907VmXuThAN1jOWTrJM25M2JMZfGols7aDqMnLjxqavMIH3ZSYiXojBvnX5EsljW
3RK7YOG7hjmWHuSlxI99yTsWvNhIQbpn0Z6YuvIcTttrpRTO+Eb5Ydfywol3fnsP
cA9ho3wviQi9VShOli4DkB1S/myEUgYT+VpVkZRUF1slSy2IpJfNTKkwghjb3M1c
eQYzkv7W/8v/rNqjjYXcOOqCjsznK4J7I15eg4FwtonwQhB+v9vA6l5OwTJxeFc/
78EA5xYhlyGIpxZpduzmnZdSZ+sSHvQOV5xGfwfFmvebiVRJJUTsbve41lAIhUzk
is0h4Vtbmj9ft8J/cV+Wt63ORYPGG+IPhldmMNme7CBqWHnlFUZcfDTiI++lTDy6
BJxtGpPjpkos6EcBYea0or96dWvlMM/f8qyQ/IWKV1udwM0b7+iBvnB45/N3s1bd
bPQ7KVdyfX1dHDXRymPAaMXe0eNMSYF2aS/+CRNxpwt+gjQbWwvMeIChXftQu1xP
Iq63ukltTkJuljVv+5w58/6NgK6bD/YOraUmlQJdYS3M+Wgj0zi02GP5RIVYdX19
OGa5KD7chqtUqEBz3uZhEKKrM2Zu4izUiS4nXhJuNCkZNQomQWcRhjr90d+JvEyt
7OWj5ivC0n0UB1tVwSq9IgUTFntkRUme7O7yg0hcjmebvROPyuRv0mJKYVIvCIQH
FNhN2t/DciodjqE6+KSZ7py6RNs/Lx+sxW1MUCmsIEzuML+eamD6JEtoEcWM6viD
lVGzRPNWpUlBqU8AcavRisCUsgcYl+z0BW6ueBcD++wapc22kbOTCfDOMyDEN2dE
tHY5Jp/mbh1DJvE96pz5lJpOKnmCAIEaKxZ+mDtmp2LR8ZiLYib4M8cQpzJbrGfl
zTwJuZuCUHGzTlMIRSAYo5Poq+It5vgRyFPFY35y1UMsp5JG0YNzMYUZI5yjIu3Y
IfPH5hF75nxn+HiVOjp3Har0hDcuPnv4zDOND3KaeJmQyOLkcH+zxjcJHQzHzNdL
G7khWH9LIDcK1PDZrgbhD0VJQL7GysD2tgfjrnws/UKOUfn2APMaTRehnXIPVVP4
4JueuLfUKJUGZee56DnVloWg2sxJuWksGanM6GlYyAP/uIB3ZfDYL8pQw13p6bbT
XG5QjyZK+4z2Z6WN856IC+rKUPloOqO2uf7XHNpBbb4TSX4lX6273ng3gTXXquP6
Il7fvy2EGcr7asks7/igt4vqYCjpZQrBOQP8IKrytMSm1S4c18rOTZ5Vj/WB/nHN
ioX2eAuz2IsQYvrlyPxAfomGzAu/J6qlyyD5m9IHhC9rnxae5QdbPaWnzq797Zdi
A/Gec8nxWVSf/N2j4one2Tqzf1R5FTT+uUfOc3JZoEjeXECBRI8JghjSR8L4saA1
pXnzDJ1b6ZySeytwDTm+YaVmzUlX7xt/HHU/8iMcE0eUIy82j1nQiBwMEif89WNC
E8HPZOZmogBhxPqmOsdEKBsAZznNW4evBt4yccN5fF0CClOP791A72al2X8Qkqky
hMPwFZKVPoCYMgTYzxlhJ7gyPOt+cT8IO0oBAh2G51YYFPQCnpcR+b6o9waLpvDi
00a+a3Z7TxFx5TTrxgfuVzzYWjYdJRoH7Bo8+LMt+szclqr9qYaiDoPll++HmQ7V
Q2jD2q0cpvQBoEr/t9pDKXJZyW1yLO8RJ5A7jvGKPqAaXFz+hdsuLl2z37Gz8uTj
pa5QAJ+EdBISPEQzvTN+LrmW5Gc4VJiudEJfsaF6fqc9G+SeILQZdUX5JUd7I1a6
ZEcaYl8QSEpysoLcczKeP6ktbq/NlFrqfynrDNFDjRBThXUOjXv7dShb8ZlKyvr2
xlGjF8+JD1PjmpPFc6JXiFBPYyXq4pw8p/7gfKmE4YQ1oYbzHyKwmJXsDE0seHnu
v+e+mZE2QHHEWHo8N4jj+2dMhLRcwpsSOftxt4cGFSo/rZxFAbTJtHi8eSf5FZTp
Hnyh8hVC4kddsuq08tN1sJJVyN7pVAbbMWFoX7AXbIND90ALgRiIkp+KeHu5DLf8
uPIcLpEvV0TE4fnb9o/oanKSs3nbefOdDrYkyXZ+Y/YCDzSqWSNKIcOh42TuMGCb
iEbdqe1ztJvDJxWL87HIsGSchPfiyo3RDntHEEdbZpm3X7ch6PP0Z1cX31Rkasv/
ayfsWqwJsUgySIzlGI+NX/XucRWItNshzFDVWTA49ko5t0BgurCzCi5cHmjGLmLp
c4m1NkATO8wGPC2s0zq4hsciec0yv7qGYT8/Pp/Usg371vrIej9Cva+qLF1O/RRl
6YTuo4MY7zimzNiykm8F3ViJ2kkt8zJiINLw1GCnbwEXz+PFm5mOWbecIGzZBEw1
lKE7XQVFHGXACFKovNSikUzlaOHM3NgJglP4raETeFDsY9luyXY8TgfOIDhVz5Z0
qdWlq3SkOWWYLC2ZEIj5ogExA2sm+E9YMNku3qUt5kyLniVlRmB8XtAL+3M74qxj
3Z2xnScA7rsoO2BHBYNFhy1wSzWLL9/MI07R1hDu7G13z6gZMsJFgYIQi0gO6qIH
2AqNhm3av2ZfyJty1RjaSbTs/Q8hzZdgQckcf2rKglvWij6DoQRoNg2dOMdAQSFA
SBAmCLb4zyYDbZ8Bepo7L5PKwFDxtumNgCRLWC2WqHM1exkDxSvtR/O2MHUeFOho
gQWqO7CMJ6OzI3o0/cATsxq0xGVn7gCZrJALA4/UFnRpAy8sPzo1tWLfz/KyeqB/
AYDIq/rq8e9WoDAG9I3yhCWGX82eybtc5HnSk9NtWDX5XsDfL8CLn8JpRoi/tXaI
HcNH543t5xJI/aRi7LMt0LFrfaQoBC333QV6gPu5CcxRHZjt4JZ9r7ag6pdgbakY
lKzRjNoZayKALU/WR3lpG/4iFuyeqmkjbeNwGi4TC3FtuD1gOy7Fh3y+ZT96hcLU
AF46446zCKUgOAkMVcHGCDWENz/aL1FePWn/bbTSeNN54bmEhtLyeZu2uX0c70VM
3Ng2WMNT9qjBVkVxt7FqOFGmKQ8v3NNZVQiWuF+KuF82yZJp+KkJJOkyM7K+dzw3
L2K4t9VMBzxPQEACLM7UV/EbGpNMAtC8CnDGIoFjM3lSaTeWt9bwXUtAwzU32tP/
ISwqmhY3+Kh3pUtf0i+nYkj+guBQZZ5h3w/2JgW9PhJNuTjN01zJX2XwTX9RNQwZ
/gkdfYxtSuOzuUNF/MkR5z5Y43i7r8Y04qppbulFEbOsamoQ099bB4wxoKYJwVQg
SFb2N8toNJ4qSFZwWoxesjOAGsEMRzgjYF0SHnDqHfnpSMsBKs7uJ0CiYJc01qCW
6oRZJuCen/TPJ//kDOTnFL7auqnS2KHN10/thhX/ZfGcdEjsipVvCoNbf/oZrkg/
1iKLfMWEeS7HPZHeu8LqKa0ccesT6Zv3bEoDlvpcu1ycYdA8sI7+BK0tq9pXgnzQ
xbNVNSQ2UBL8JwkaoetjEKzwVpieDUzyEKK+wLLdhobSA8eIEJBrKTpfkZ8M/BP4
ZD1S2QQ4y8near6UteGI7i/dwb8fP7QR5EO/EUSanpf0YJjqB3EITdDJE+FV3/w0
4LA4V1GKr0q5LI1nsD5a7EB8SileRVZKB0PFUo7dxWALhp38rZHxeECcwHw/pV7x
3AzIq8Q1Aw3Gnv/4Kgpy1vJU6ZJAovbn9V0j0/Ivvxr6AY7AGlr4c2vGCnUT728d
KlixROe3HxiKJ/M5Nt8p8EsVGry1Pv0ALzYpybHq5WOGfjJobSjsF8d7kPqDb+8d
afZru6xS2c3acZyun5ACfZ/zn1qYEF8gmlyyQ6fKy1ayrijz5NWi0hqOqwMT/c7g
h6xhNO4pa4vxfHoAXrpBJsAhq5Y9sdXIAQZZsrmkUnds3DkOkdxq+1hRgH3BQHEm
9NccK4BnN4FWhKJUpm82gKa2CUYf0VMScZZjK4cMAT79avmaDYfqOSHDXgZ84xDH
ODjw7YC2PxsvK6qnU4fAGlxZHAfCfT4i8P0fG52McxZLUwcLZdtbjEqeHPWbbBfy
H5xJ8zUgbnqO9E1CF7hJrdErwiEYt8iNgz5NVsko7IcYF6RftN4AsDI7L2C9TeQN
tx3/w+pM4zP8NhPF5uApXgcN+QkBQWJEkdRFFsqnICgpwxbnV6Y0sLtcOPU7NtCW
R6k9zgPR2gg+SnmfaZ7FGADun7SU0+5+xl/5XGjCcVar30SwREiay8uEZJxMw92Z
E8sUU2mXUzTGPqA5WstwPHDh8SDAhAZeDs3vl4R5nKpk7pBoHpX4FYx3fuZw3h2C
gjVvMNFiuYPPwoZFBYU+/l5oodGStZRZX5FkWGWQgYaXZLDRvhEPsVgKQGccwyd1
e/pLyshlQGGlqMy9Swy4QvrFIInXMTlx2H9JgbO7W+QLNusj6fatriMzPVjKLqi3
5J5k1UbcrEhveYKB4pqy/zWe9BIvJYxj2KWqMRx2xD14wwMPc4QiEsSEhWlD8+NE
NefySl+D+Zxs0yRsbtPE/B3d5F55GIDz/jT32i4ciUTgkmwFDoA2QvFpSysir/Me
mgHlM9t4i8ley8b8lcgtnwGY7hjnPv2NF5V2ej4uBH+9oWsWvULA7q/jaFiasBva
QKBjc3Zb+1jaoRuNoQgEo13CTsuBnGb6PjqhO326hn2fSVQZ6M81VpasjGg1MBZh
Ez91lf6q8vFShp6OOJPENc76Q3XeKjeJWbCFkcmweXooARqq/hAyogHsjkx+HkBg
5OMrc3LEzw9zX2/vP+6dygr4XbZP4gIo8sR3yfg3yW8QcjGYlA9MwKqALEASEuEx
PQuoI/99Tpaq3GK8S14DMjwJukeo6f5GG8UHyj7Gzky/OuO9oRyOeSoRImdkHj3V
RRpbOZtAWtYR+GOAg/1/fKZ4PbKFzmGrpELW7Vb+UTsQ9xdGJfeIupGt+q32He1u
HhJ/tskb9hFlUmvaPyceEGkfnPsBIgNqmAbytMr/7GoXUnmhzOqUVtKe2YkFAVPS
Lhy8jPM0xM2HMkznH9bzOxLJNxCdG4U5tY0vcVuLPHr39rVfdZwVsJEPj9pENW5B
EAS6H9mwMoVaN/aYo8LwgOzEEvUh97ZcWevAvJIaQ5bsdqeu+fNAIF5DTJCENwyc
modoMx0wjfVT9U9Qmq66+XiUB4aa4/h6iPTmUHthuozNfR09a2hc/2fYKHc4Rkuq
qa15nygtK/Xv+ZwWPtJ3j6v4PYwKjJ0xmeQrQMwF2q6LFsu4tFtfbz5X3XGjFFt6
nfU5bQOp2UD4fE+IMgoOhLcppwmAad5U9fivy4kfU0eco2CwXXtBRdt+QVGmyS5b
0eACrUxGrDmgW4ZZGCBv52MYIRqn8t9VVifzRpjupiZPSKB+EhjYoPSsXi5TVBJC
uSnubymzwDzIpT2x3ZHfFHImdLGbCx4Xa6oB1I4mSAhXtuZqIpvhziN5g6s7MfD2
aZWtHXwIRcNr4rHwVzMKCwbsu8bgyfzgHG9WaHqmbW/nkwLnFmZYIh7iHCbxaFsa
aRy84b6RUC3jz/Liq8iq/uY/r0Yv0fNBDJAaMgWP5QU8RYCs/LTECAZb+Brcv221
ZyYAWq6nL/JfGcNdcCEDexON+ZJTUDpF+OYilka/uj1C968DpH2fsEEsZeNiJdAB
dxoMBSzLzheVWLtdfH/roWXSKKC5wJlykaJyaQwYobEDCe62BQEreo0gG67Vzjpx
BwPecvOQaBzVzPIidgLR0WP+dn4xm4V/KDyPBM05VRmjWURO2MluvHg40PE7Uw39
8Wj3ZJuwEuoGxVP6ECQqH2/oaWJJ9JieEczGIy1jwBSbzWH+EjHFr+micawA+AcH
HVdx8crMuwZjujYdgPKNwk3whT+vnIVywcoknn040KqAW4QskrlqdARQkD2Xi+eK
J5cZnbuyR+TkwDKFYWkDaw5ACs6pcGJSKtRBmjUHs4ojIUNKKuJqeX9hJa2W/54f
pC7YIRx+D2MvGAY5nk1wOpv+DuADUUgq6G7kPNMFo8CLDqND//Ad8bsFVhpgOc7t
m6nf4UMWb29bRwXi9aXpMzFADVPFhgVdeA8nTYQMtOVphKn3r+jEiOacsZ7f9ECy
S9BzgEUoCXQVA6k2ndryHug8ep8NddNgpEdmb/QaTZJXhvgu8qB39YnOyj2PZwId
FpfMXcSAfC9XSdgs3kbIXpAZLU7vcPQGsb4bQjvY1lukRyAv1w+0mj/IBigwu3iG
UtGza1II8Vx+nlFuewZWmdAO28NMr0N15/VzIhD71r4s/gKWoSgTxhdSN8NvlIzn
C6h5MlrV0CGmgvuJ2+WU1ep/ouUzNWO48S8cdjS+VL1T+tnrrMH4PCsDzYgBRwyE
+/vpvtNcVkWhxz1in7qG68nXXRKQ7pLCJhZ/zEmArwy2fX2ZH2l7Y/4UjySFHvWQ
rZjzVStinwVN0xYaLreSAhS2/WSpb8ZcWaXL0CtXaMXGAhU6+hEd+UHykVwhrP7E
Mces27A8SrvtFpUq+GjBIfAuvt8bLU6vb6IWfGnoHnz9aM67oeKMGAhSnstS8sH3
s1bdS7DYMP3eMSFVTRhgp8VkpHyJz5St3TRxXWrCO3+iACgLKTQfd4FZOkU65+4K
BPu8+sO0JX3n6T8VtMEM7TNtiWjnpBizW/IpMS4Vx8ccQ3Qw09VBDke49FTDtIJ+
G9pCKRbIc726sZMwfPmfJIt31s925BQPByESAwiOAS+dGlsNmOlorVBcE5kwEY6Z
b3HEaUyW8HxTyhf1U3+eP3jNLkZBDmovMn04ktScF74OTjsqAVjSKBJnLBYBKLdS
BWTmD4A3bMPuhQywon1fPRaJPNrz6SX+6tOwTA8xOf97W463Qf+R7bUTJSpN63cR
e3md6SxU1FzXtjW+yQzRodCJmpAmic6tfB71zR+Cje10Hv4C16SqRX9XdVq9dGTD
9Yhi3v9uMJciOdqJzVrHopS8WLivY5ozPtGn1lfmuXykmX7eVelQTwau8+TZUV+u
QUS6K/l3u9xfymc/fbTAXxIprduD3fjrNwtySgAz8Oy0vuWqaBOLskuk82HPVcSD
kVrHkBVzwSky0A6avhC28Q2AgjRhq4ydvhDc3HFCy0cSz0HRKLPOxLv5GfvTVnB/
/Qa5Chpta4vnic9V8la/rGxdJ7bVVV0RdrPLCXNaFwNviK7k74uXMRdqjPXeCVkZ
wbvTww1txHgWvO3aI0oBEx3zVOTSR6oaNsXDIxWIOpAyk+eacRFMzFM+1CKhakPx
Y2n3Fo4S3ZfePRZ98qxE1+yFnQEtRtVjzciCF3kyTdP7LMXGUYXodxOAjotpON9Q
RBtnYsMxKueFnZJAawcQ8WiVPGG47gPDJqsenhfFXV270Nkl/rVTidr5DbrNiiei
XO/ajJcTisUeLeJz0hwSDE0gTLieeiH+8x+7MyoTc59e65xmlMIOEvSa/eQ4XY6F
7p1vlMPC0AiGlmsSDjrjm3TONhxWbrsSozu9zo+CF9dcZindrsdH57ADPnYVULz8
Uhqt+0cL0dog6isoC2KMUBcLsG8kpE2INO7H0hD5hv3ooWgNmwym+5G1LYifKp7d
rRI6qfUZZQJJD+rAuFrTNWwSiyzTjyjrJ/PNpd5VcL+LclQUtPE5JPn9PTOy7d9u
iVnKuwntKV22BkVnRyIJ+iH+7NQ25rA+zH7uEbbsmSU03wi6eqwr8xj475OsYNuU
bH+xYQLc39EufCYK7NHeg+hRgs2EANu4OSfhwV/5GoJyneDE44lSAMyqJnMQviMS
CA8OxQPbn6ALCeaSSNIUijCFDosaWtaHjdvoDKD73IpVYxdSW2s8wMJzhNRTeW7F
707xGWpGqzlX6B7ksCm9sI32QfChojLmh0nTGnqU3SZQloTJhLpQqkhfHn/PkfwU
Bhsnp3xHmdnwIlZvOruTY+wh6Cj4T8zoCA8gV6OO+BRI/ajC2FjuICIgJotw5uV5
XhduskmibzIyh3jQAeKlK1GTdsi3yx5wIu7Ha5zmK0W53J/61OEWFmGzBHRQj5Cu
UI5hEmo8V0K77C36xToPO8IBUOsh2iWfeyH1r2IGdhz/hvWdB1cIDU/Z+Cz3EbbD
ucA8c6qtk6IsTnRKhmPmd2KM8cg68pfLzwXaSjDL/aJQ/TKTZQ+hR/BFOj5Y6W8+
HDSn+IMDwzVrP+PazrA25AnYZOtT9Yvy8Z/SlV1SNjef09NFNVv50BID7Sd2BfeF
Ln7RS77kcKwg5C+tQP0bbkn0cK02Q+s67IjFhwdks6rm/uoAJw5H/FzKNVM61u0w
UJrA2pwZmC9tD7DPOpslTc6sGN8EEdkQNNhteUKC49aclEWyVTwSvxzt/4FQZryz
Ayg40oh1PNRZkT/NBj3OF33fj4G+aS+WE9tT86cejv4Tam/sWCW7LQjDfMTYeLq8
We2ewxUlWEjc+2gdIBNM49UFPrvvrw83/EHrEt+xHzGKQZlU11wUvphRQZVlBtPC
jxA4VVzHRTwiYWj6x8+SYd0L0J4Y0j73iEFVrqEetkpApzdnxXNILKPQtd4qTCSt
jlJZ3z7h44UGwW5AnCZS50GDZdmqYwBhr4VHayqkEa8b1LXsOwDXISf3bbqiC3yF
N4d08LoI4caL9PjdwatKbApS3t/hC/GOaAwhVHkT2czYkOAc7KXJVFyO3gFOFi7x
j1iZMcrvuRHrl9w45bT4MEfHPNGuDAmZWJGXjrKXXpHUSkJN3ylk9bi3iCqKcJMj
To0n5m5OAgwQjzqLbeG7In35JepQ0IRgrrj/Imh4nEoTfIuHSryxEL/lSW5ttot6
HjorFlaB4lJCkpGJIKpsBHln7t0rrtG26Fpt61vav5Rko6euyjDFGeeqAK4K4H3k
WXIda4eu/LQOULnLrrcnpcXxM/gzZBylpmxBH4kUbEVCd1ECLbk4UPZpiv1mER81
5yivdc5l+Apg0/Ed484YEXvJunTqESE1smoBOv64g376Cs53iTkGZFBV7sLOnkJc
AaUoab3gBvjHYa9yo4PDbanfied4GiUXRObX+ExUC0CHEzfsQG3jWLb1wI/2l4Lr
WAqyJUqfz3zsq3tXUPgwYVTrY6IVY7G4De1G/kqBZ1CmJgtDkRpO6iGBhpBQ6GH+
Ggt90Sy1M5UCkhLmZA/shBrJLWGeEZkfCNUniOQs3uNSm72uWrvovrYstzzpVNHd
WH2XiBHQsr84Nriwv+/WoEUKLiONN/WXDhUGjyfXewb1FnlSywvUIM6rAb08fNKr
RWqEiiXHML0/Wfnwi761sjb1ehgZoLVXhbpE/HYSMKBH+eDWXmLN2ybR5lAMXkWM
Cb5zOOa/rT3wd/sGcdGQR4PcI8KIbA7Ql/lCmWPaqFB6f2Cb+Y+nUNFmzSrPm/ge
LepxcT2Bel1YeuklHJAXp9flUZK2X7TBrfBES/9VNuwbsSo6ZEwYgkxX+IJjUap2
oSZrId6y623WIMaOG28Bs9c0SQiaOruq3B9fD7G8CEYIrZOrJ1pqr7mUiwCKAS35
PpmM43VBBxhB9L6biViRxiYTqFcQb/HQx/r6DxEr14SSJOt/RL1QNyu3I/ZcDPox
cVcMGkvOtdB4NLAYHates7XcfY2ibuYPUzs0w5RWll6N8oPZ4TSKa26Jmdp9UrZY
LLmEcP0qkZMD92U3maF5jKHCoQOk6DAhz4OL8mgJpjqldifi32tPvqG0UrF0XCjc
dAaK9XyGXVBCIdO9rrs6r3Zefug6GE87NzZeqv2V6lOl2GC0nDkpj9EvaNcWxECG
9oMFfCfK2Co2UbvPAYM5FsLcdTR8Umiyon75Ivf91pDzDcgocq66h8CfHj2Gpn1v
OwVku3ng5FXS88JWD8Oo1VIMT0jYuBBZIepvCE4Pk3q8DN+PD52hWOZGjiahPFsp
JOvjysn33q+s6B8RUg+3SeNM/hSERGjTL7BlPT5N402h9F9zYsQodTmr7XIARMvi
Q+ZmWIggstYUEr766yzKyX8aj71mkKnb7jJkjM1gYms38bohxBhM4WT83dr/pG4Z
YHeo6lSTHM1FpqTq0Ug+Km0rwsfL+4Cy7K9anooP8rGlFPSfEV+in/aJzBYI0dIN
IVDNAEYFVRBFy2EGxZZKW2YWdYHmonV0Mk7+aevqybHBzBpn9mHVXyYVtTV92pDQ
Y61kZ9wgG2EsrlMEeCJJih4F7kJwisD0N1FuAwBmkHY01DU9NXWMfZks3uBCIf7X
7V4qn2dZRGM3pLpUeLMfbYhzlWJ2KY+CXIdKWXE01sESuhTvvSIZ1+g2UuCn23f5
ZGTFUI2O0CgeXg7wRUoO1DufpyNbPTgcdMyWyibiWO0wUieme6xuptyh8gQcYHCq
WyE8KplpqXKx7W4CALijr+fLA1Yy3ckIzo0d1Qrmy0v6KLfCkJ7AB9MtKbFE1OwD
NXhPTqLpADoj2NkpqKS27/vvNBfZqMp0lSyA4ETAkjyHXZnzGOdwUeoleIJEVsQy
U5GWfiisMcS3A+a1ZSdtUw+Hy4N18i95l6QhgyZHhVNvFwoePcTOKaFcAyUSLaCC
6buBxgpXeFQJFEanTlKQyt+ow92mcMENssRaXuaRMO4qzVxnxq4ezRJQvQGx46+E
rWlDAbswPyfK4Sntko6eBPOr2V5/YetD/QxCRxMobQuOVDGPvDZ1SFwYTiTx6GQ7
Z05m71CXigH2DpPBaGQBB7bNkoVhzItfFSTujEeCGIXJ4p/EQaitu7bsOrwRG59Z
2RtOK0FDvSXqbbPGTAEagQBaWFJQBEqtrlfAaXa+Q7olUkPPRWc4bOMxy9pQuv1Q
luIsOhuMOEwRY6nyw1WR+ZeJTVaCzVOZhOwIezw3YN524y16nBA+ONnDRJH/4S0T
Ww7eif5aNBzE5bL/kYRSK+CVU0P4c0xKMH5YCMaL4ZkDFS8Oq5YovaDpTqwg58Xs
bkwhEg9XHV+2PU9r+422qBz+ikl6vZ/zZD4yR+CZxvbE0WKHI9RoJMUONfXMfbQR
UzpWaZgZhbuxNGm054EEVlnfkPDSb6AKEzrBm5BcshdC2bcnawiq9tyQRoWMjTbV
Q3uOHmvzGtb3yJP5unBUsyQrkFeY96xDfhle1Z0WZYMNFfivrlNbm1AlBvqDGGk6
E3zs5tdP/nKx/XqrqU8zOpthz5Y32a3joW2VGfm0HwzGZhQP7jpMHkg85HDHk2QW
srPR/ljNgWDVdgyAXkLnOZDpvNxarfLHv1m2KYYzfqiaDsK51Z7Nn++Scvu5kZcS
lWWXkIHx8FYTD1kvn/3UgqXf3400wNuFeRAC//NO5yAAK592mXlW9FwQ2rzug7BE
Cye4SOdZCSRK08Bcomd1IQlnU3o8bxPVzw7uvhwiEL/mEX4f27mm/DS8vUJL5JRd
nstZ6jFeF1cFvCsJFLWDHwc6N2Nk69OLICICSqnDP8zOf10M+yZkMsQIelSEljpb
9JxbN+yS2S0iSPpGoSsAEt+LLS6QLcOvqcI+rCKgVfMet7/XND9RyuyVvFquMB0t
wvoIC0Bxe2zWPnY1eQT2mm14jNuySPZy325iNEgR1K3JJpRJ2XKULv8kRxtq/wov
RfXMtWFqroz6ucpdtRiMk1eceUAcevETit6sxaGoOl/C3MaP/BfYYAAUnHxY3G9A
WVu5LswYHH0FnkFgaqepFtLUdQ/3JPbw8Jq4Sn7VmWuzPG3AoY43Php07Yfa8BLl
ZTngJsx6/FPOa5vZD45nf2tMeK8A9NqohdPR9Dkx/pj8c8IWXORkvYuTTy+8H1lb
rbfYb6d2R2RS00ZYDQcrVQvovYVggdmvHxbmkwZq9E8tDT7PeO1n+qlSTBVVAxd8
cwzLB9xUOxlimc9jzjgHHjQfkXEAo16aTuH9DBO0pB9MaRtgX1InrTPNopgSh/Fq
a22ZaPbk69VQYyf7wTgn2aABfNqkYU/UMcpsRiFjPs2NWTnQbHadckhp1UD7920Q
He9Z8AMyU6JqvF5rMfEXCCLnMJhE/aAiy3SAe7T6Clz/5eFt3VlT0/nTfoEF4tAu
1f+hgR79ci8igXMx6y8VWl0xuVeAxX/pKbhEiIIkRKn1lW1NZD7a0k4q3G2ZzHa6
LxqxbV8hdrsI6oglVQZ3B29Ou/Thh8QBxEpL/d3BREqk3dpthu1lqHWdHsuiQFqm
QJWdF22M8nOnFgBfa2M6peSZxd/z/Q5MQUFrIVdORmUKpExbA4vW1Uttq8NtEikt
KDxXfVaUvPnYYp3iZ9LZ1+95RdfsRm6HI7qzkeDVIjvPdN2+Zs2tQjyjBPkfn7DM
W4hLAZ+eOWpg5Cv6nx60P//BKQ17+YuiFALC2U7xmKamn3nlWAyc26XcjOicncmP
tImykkfhFuEtSP/xdIu58GtQDvQyC2YcThnIKmfW3BedDsnSrGxVXX0zXfH8Eic3
lULDaMtL4NQQrP7q2SFvGLzP76x6CLLqTaHQkd1iELbKrErOPg7y5P86t5OcPA6Y
YgilN93RNAO3OZLhbUo7tZtThbj/AzH8BZbhwhGt0rTGTMQ2a7KKxQsOI6bK0Xvm
aZfJUG4h1RwBB2gXKnhX8KM3wa/Ue1K//FXmzh4l997Z8UGmjBpkt+lEY6Bw0RNT
m41pBO7SnPjqrnaJquDONF2hXsA/Yubxk74FgHRUnSusqkP6cAG/c0EEd9CZXhQ1
YheurDFgZztS67m+ltmC3TQjmALvNjJfLyQVQ9mM8hF3KAb1xtpmK1C1RtIefXkE
Dxxrysn6cCutR0KZ4csXSV/hOSSjl8Mul+BEpxvOaG9XJWnwCTD+05RuomKAw0Jo
ZLnypHy1HvDJsCUTI9/pTYHRiTNA28ygtINP+Qk85imgounWIY3hV2sUov2h0yAi
noWTKLnaPp9rOCLwbJwRBf6KSu6VIqMBfWIi7lXaf8QxwRT27tSVREXUjkU/dHLC
cjaO7c7WLgB4TJ8Megh4DuxwERt4GZ8GoS48roLU5RW40YM9g3B/szvTQzZ76MlM
uL3XF+x2tsUPJgdqhishGfQuUJ5XRmwSs9wKZuIHm4RNUlnUdVyhwJzCssrry97i
ijogSPMdrv260ezRvI1K1uQ6G/FJnoogBoCrgRj96DmGn09vOI9BGpv1midwnM3M
QfRX/xkT0Qj+dTqMW0j3sVFukLdVU64R6aSWNk4Qkz/9SfWIKPt7rJLTYul+wWGJ
D6FVAxDmvk+7KkWeaubxqv7l93jIE56LIkY7d8S1DDTAUlw2PcWli0pD8coURXjK
AFJ5EQbOl09Yq7zNWa5GURMJ1opHAl1BvzqM3oQWQesobQgPHVWdqD9Mzbi7yBzG
MUAkJGuTTeCQm9wrxS5h+hKdNrdftsmf4yE4hMqJvYjdomQ0Jl0riaN5IRZf2+eT
9ZMcoWdrSUkn6Nl1AQdx3kT4GT8xtPf/VHZ+8EkSLrNlN/8MEO5EmSQg1MOoJgnb
jt83jzRipIxtaRAYGE0WVAUgB9p8kKkld7FLdtTfY9HdFwRLgJvUoz0Wqr3hznO8
ZtKWKt83yVuQNKCPKDnTLCL/I0sk6CjrUeP0OLT62AHHCQd+3+Lk4SmQLgVQitFW
OKIx3XsROejbF1vxIFFqPFpItbg+c++New7xfLjnFSOyQmTCIVIob6yopJXLKsUH
6/n8DvXd76ET38yapf0Mhz6nBQr9Cmb1mE3l+9NQUkKF9KL7VQ4GxLpeFAWxRwO7
j3FkTpj79KCFvcEiXpP2F4EtbVXj1EfsztLXcK5PiJx5m1Df00cGr1gDQPLkoZco
uxo3lzDubFRnr/3fDyuq09qQuCckI386d8x3zDMe3io7TeIeReVJ17GBWiM3w00e
XXhyr/JGPaAyyUwq43K966HNdNOt9mGwGU3xS4PTX09uTOtcnAgOIJW95eB7FhaK
ZZRIT20powF6g8OmXWlKPK/9MKycRXm6OEy4+Xo4PRvqqQDhp5fZu9guiAempyW9
aP15FprW8iSyFTCgm7u94TaUPRxJnZQgSdOAmfGFm1harGDa+0zUCtL081Ddhfuw
zgWnV+hrWeRUeKC3QaIPKDSfC75mFwrpBFkxk2pPA+oNYlTrlktzx4PKZkQiC8BW
Y8XVhM3BrIP+JZiop4s7D2HS+NnQw4pBJyoJvtIGJQcVJwFrVQ4Bw13Y1VsEzFtn
X9Jj+Y0qZ/A3s6ArgyxHgBngN7PCyzHrzp1KL9yugLM6Wl+YIfM0fbA/JTTjqi2D
EPk7NHwOvxHeJjaiEvJmBHL8VZTdAasq13tw2x+eFaXdiUOri8dt1h4ywIc9VC3K
0tfGBiqU1JX2TH5ZL7LeZys+at7Scgo6tg53PNbiOtpPZzeI77UYDPguJVSiY/Pi
ztRN3atS6iV02mIkFx1UphaCWp6aopQF4Tn8S0w/eechQ/jV5U9kHET9jBhO+wH5
dRRmP5fOV7rYFwoP9DmDVTq4G5gr/xaHbT4OIauKpmXtahi2AZSZyeWuHVJIHheP
4f4mU0BzMTV5gieHaq8ku1nSGzBo8wv8Oy2iypdlPI6LhhFyDF4pMtoY1c28wkfx
MxxLbSv5fJZDL36RZFKVW9M4NDU9cNK9fhOBoR68UAnmHBsmIUMMuyeMelSt2dtL
pKKkP0NNkBKd5rwlcu+egNZk+2fE5tXNRNyc7IPryIJ3jvTG+uHC5/wy2FTvPh+T
eRa46Zi9Ij7dxuAh1lFQj+t27RYXdYGpP0aWTz9aOczRvn9vuPU9l2yeIvuYEwVB
aLt/rm86qSgJJIdLL5aH/t355Dw/FiqJv4qB4GjfRBdJzCHubdy8tE75egU5Sfcy
+fXTJPjBZ3PhXF3GAw7n6q0PXUbqldH21XfhsDPIIwLFGBSzh4s5ZGH5w+A8ZxdC
gDW1zWONJ2KAWbUvo1crEyPKSppPIZ3H0QdNMX9zatGCxQ0yoF5Sr44Tak1T652i
o6VWpcWcCZmzb3sR88EcLJVjGEH5lgSrUItfTfvpPjXb8IW97QS7kp2s+B77+Koh
i3vMspgvPvGlAsR531ve703x67zYWzyCSCojiguAjJwZ/qFp+TaUAqa5bVoj8qee
qPdK8xhP3GfHHsJ5VqAUlVcAbdbQAUxTdRT29KVi20l2dWpJJRmzVZx+awEkjI0a
7uu0eg1xkFQPVywc0TYeEEAUrCZb4GumA+NXg5TQm3bSdPR7SXMCPeHJwJ76omsr
j1jcZ1DYDgq7YKEfunn4X9k0pVdVruwCNxQ4W89dDs3Ft3x60KDva3tGOFGpGiq2
pBhvXjbFzJzHfBLVTLeRxrLXLUl8Q/3rAmKBqgUWmEEcrlo/Ib/4avubCw2c3ItX
pBIsP3SCgoqHuJY2HqGPG/0tE12OjGPzFcmqcL0C63ILla4hznxi7dmcWzp1itee
Csu+b6lOy+43uLideAs46khwVDjqPWXksLYOXxFpVcBvYGXw86k44Q06pfGRDfcx
hxkdwmHHdxbFff498qiEMX22A6VBNv7JvxqVF35uk7FApwHW+ynUp9sueISx0+9y
5ftT+HHn+wOuVwwbqFaSFS2SHLVT2NaEe/xO0gA/wOMgBsiaN4YOkMAKKB2DReqA
aYTZLrM2H6DmG3MmZbBYEEP38/04613GkCJqeO4Krry3BKpnMSwmJj7DYQEN9BFI
ROkvnzim6v9GMiZ86b3e3NhDP7wLxc2Y91raJMWsMoAeZyx/DsN3AeAFBomP54Fg
c1eFV/YioWnbChF4Lm5VPQSEbYl7pPbGNdxYkgZ/ZyvZnE3DNd80aeO+lj4Y0/ah
jYm3Tf7Tj1tMz03peIOPbmmlknk1YQrdiAH0lOQ37M+nibKxgtCUgMEMgRSnUOia
ejyfDrYhbLJ25UT3Hm8EHb61o0UVP+euBXfcOQl1lszI22fZIQ97Kg1mQzCQU+aA
C2HVpZAAeQjzEV5rFC5G4HG1Ea4NTdKdixAk1Q8oN3yJHmnoaDyJ4XgasihMdJnW
5oO9JkAOERvp6Kq4TJ4ii88iMV0hQBr/EbLhNkZFnHlNQK9Q6fHvqWiAAXXI8neb
cBDG5Eg+/ByDBq5F3/qIi/aI/Y4bNbk6LONvO5XvjOjupRwz1HXhwHRy4EpGSHB1
5RAcLw6wb73lFqaIo1SEf/L7/ymp2k/Y+0cxLw+7SpvDjFcmKVL47i2MigsZbAXR
9BI/7tnCJXNNWvrvYiBO1jCGYjB3EyOxKQ3pl7kD0SPj8bXsERmEEyiDQVaP/IdK
HTmflgo4tZMXejYDwjrqyB/IifVGuU/l3FrFJFCWBePW6bagrUwyt8GVVxWUv98k
ond+J6cg77mhbWU60r1t1o+mgOXHGZnqH6fGBw5RNPVMc2BXGKnqa9ajU64TT7qf
/ZnNUrlPKFmhXfAN53XadRwUYrlthjW8em/QBZ0Amq6uHLioQ/zqaLFGNUrAjG/Z
+sbmAc24G8J+8GseWYtgUBf9U9+gm6x4Mma8fNTmAcqFYtVBVBfP79iJ7Pa1J5yZ
iZnhrAwssIClVMO3HxCIipVJF0f8Wk0hPR3oOBHGOSAPCLe8UAXhuIVherwRdrCW
I5I7rEmcJ1dZVYN27X8qb3UYORiZIOw8CeYpHjUDgoE1ktjKaBXu8J71id5uIdp8
PkVVSdIdTtSLJXG/ViREwNXOmhxfBmFtte0MBLWETnLsqXLu2ZfydlpqCS1rL4rS
o3p10+W7d0bBu7Q6VjegkE6R4HtGHGbI+s7mOrx5rXz8kuNTb5V5ooLPTHxBCnk7
ZfwKgNwISwXY7jM96LYY2lt9vlHQQdMqIVECWVhC0dWwcg7DBVXPuKRkZXxwDatr
yKn/sZOsv+JFhJrxuWMdCFq6kNAE2YMFkS+7j+1kf7DrLAAO4mJW5MpF2q/ZGPOn
/GSVceGjFvTXxXC6Yvb9NCsLokOZAgWk3hqSxqFu6Yxmv8t3ZTZLMVo3PLj/vC3n
sHm/x8zH+IfuoOKx7V7YXNq2OPDTseDg3qvKoYEbJcsBFK1Xdh5RTR94uht0gkWv
0gwMwNmgX+T2D7jCcE4VZbo7j0eHGtSxXoThVCM8H/WY5XWFGxZYBAOhwrQceU5c
YhXw0oz168e3Z0LT+VcDS73gZjYrhGoFdUR2QezgLHFgD8UdMmP/FFP0Nzfh75vO
tvU59Zgxceo8oHV72uWi59/lXtCDBrJPQPpiajWWqY1kwLMrPQc2JDsPNm73IzVW
3bC4GscmSJ9ZAg0r30/ZCIXpe2XGU0HFlXCUT8ApKrP6ZwR7sLQrUUBqCFLPyuqa
b/v+ktLecKqXlAVOZ/u4/yd5RfN9S2LmsEjk1t1YZ2LwKrILoJ+oUQ1SK+y1XTs8
syuXRBBChqfNigstI3KCDT2xhafAyPcoNZlglDFBjg5+6XPD+XvRsS9O2bfOFnXi
YrP3k5tYpEOodMfJ3ayycAWZvM2O+HF6TRcrsh9J4wH26m1O1fxRdq51ps79zusZ
8yxnj+GzgVjkrSrtZWIhmXHk90srfvPHqvfR9TIq5ecCjZaa3rhtVYiigFSHL0aU
Iz1IlZW6KyS5T/Swd6N9QRHNKFTwOw0FCRH0EahxKa04ASYQjTlJA8ql81qQwlm0
A0IJtdgy1Hx3tJLnbOpFF4oOdKfR2OSZskPw54zWuN7MEdek0BQIuQ1USLT+SXgl
7gZoe+jbBkOzqHAJETyGdxkjS128QAUWx8uXvRvvjzeN5O5mwhsA7h7vMrVl4NN2
gNRKYhZ83sePI5BcD/wobfElc3FRYzdhjg/E1Qq0qSo38QeeucMZC7uqtB0V5yla
8+4YFwgfx9ZPUTBOyLkd33cNj1sYJocGQ4nCj3ZiML3DNorKEyPTKF1bASSpwBuA
YuiUXkOvSFIwPH0vwChVwVUYeuSCA2scFn+YxkVwYq5A61otMuonGvQOBgDTHcqY
X5XW2JQiDJpjjsIL+KrHg+resVN2rbp4IAUhbt2epGzsFvgHj8NhRR+oIp5xGOVN
+mK4DrJn9zjofGN3ZVYkHchoA14ZIecNJSMPX4VANT62Zt+D7nIEzANh5YvcV+yi
02/vBiGFOXWPpE7xKchOTs+yxGL08++WC51oo5fOacu34nseDuOsy5j+EkIpXTBf
2Bvllae2PQSG8vhsMKQCcPKWg9SDzOsJ7T8e75u9UmPpE+gGWBZ/fzFI0bCKcbpS
LxpjQ7mBAsTkfhA+KRmsHgQUe5/yE1EKPRvYA9qo5r4eMrD3+4YxQ8UnENhQcxwU
W1L6IFFZAsxZ8PO2cEcuTxpUtjCg69uM4nR9sK2+8rWHNixpki7AxaI99RYMjiKn
NIc35Mko6yhwqw7d7GW7P/gaXl9u1Ffd+k6fDB4k88BqcK+tZfhYCGp+CEJaPtW6
n9NU45yGeJwqoNBRUwF/d7KhZP4UrZjOm/Q6vEICy3GOExZY6DcJG2tKKOoJLr4K
1OMKdzO1z7WTg+D2x5qRqgjY4TUEtb5rmRbKAk9B8aHWYTZIlBmfeTaKCd59BM0V
RzfnxCN9qgY2KFsqG806MNeH55nYXJsH04Kpyb5UY1EeIEsb8155uYxpolis5ZPH
bXkw3cjWqwzDg2Y0MHHmqDe2Udzt7pqHzV3P2vMLMhWRsq2UwLE+pLSzlzOBjy+M
n+LbKoOksSo65S6WeuRDEqaKuFHvi2VARoKit6R8lQRBxJ8WWghYwfOVNluwGObX
x1Sli/WC7S7CbBkkAH+fA6bPRFy9qf9IKVOGKD5N/2Gcqw5Z8yGVoU84b2cjbdt9
HmmNGeq7rxZT9sGqGtL2XO6c6WMTBVOpqp1FUiuMOtSByivB+u6OvZnWYzDzIS28
A7MNQbKdfbnsfdMneC44HSE448caPrBhPzFwndM2MXzsRrpTX3Yi3kR0PG3sWMTY
Tus5NYSHoO/M7gOv+/h7qR/n/ht/eqK1xnTP1c0y37Lp2yyG2lrSAEbwxlAHRDQm
aOLzXafKE7gGc6NGxt3TKndJq7e3trM1VFh9mvxBll00vBKChDfzpxef0gxsbBmy
kl7HHAruasQjbnmdnGl6ppWN9y8bl6OVwgjy4klhCP+T9aPCBQ9vN/Fnmd2FeA3I
F0yksPkLlJewWn7i9Vhi7HAXmjnp2sJc9haWg5+awDBFm2lMlFXpgQBFz76FZoD8
XE5JhdWRDnEthQIUfdsYkpTCm7aH9R/L7fcDWW3mVeGUR6gcn4ZGz2Ik0P65DNyS
8WQwcpXsEYBZRFhzJsq9to1VokZ4j++vf7DMdZbvwDXqARTzHq1CpLrPt0PFl93K
BUOetcLmA/dPcIKFJff/St2z3MNaoNuH67Yxtwlh/vwra9dKEf8s+C/zVFZFLLOz
C8jWiI4l0peh5cRe5zb/8ijK84OdPDHYxtU2M4YYx4flDJDCfi3W14BkzhJyUgs8
FJ5EQRODNgYObAm+CIlJtGVWeUG8Gebhv8psX5XaMLUV0ePcOXlnCVP+blYfzDB8
yx/6B5o2ZtxCoT8D58JFTIPaeIZVl+JWQVkgKQ2bCDoFCSXW3VEeakCthsEfFlzP
7zUewO8KeoSGBakx0HO0VUt3fdIzAzu3TswVLhvwDOFfefZZ0NorwTJrqMMNYncc
0B0xODOgLRM7jP2srjEphgZ743rZsSRYLEhV7GHCV57xmXoHFYqSLMy2Nw2upLU6
0P30e5u7UcSzPFfz3MqKnY9A/9BqfTfcGbN/YA1mDt3mTYg5FOLhAGYkGgP+uhF8
Tsaurcq4q6aP/H95gLSZOWqsJ1PdnSWai6YElrd8JU0usDZMiCWLLuztQPkzuQSS
cEs9BEqepfBiTDxg9UQo+vHmmCbwVbXkEjzK/uIivDfYSiMCHnKDef8PD9nAqWn5
d8+Dvd7Y8t3IHT+AwMnqqLKhVHXwVXf3BaRhwRILsTYdLxUDUh2sBhtqvNWzBHjl
ifClsuwIi0R9IQkOIVfoKQ9QsDM1KXYnnJhTcwIMhPrMRpaSIeKh8ml3Hkp2Vr0d
4+wxNoivOzPD7JPkM3NrrwowmDxvDrhtDmU0Wd/1PxXzcmVs+TenCl8FzKRfsHZa
nAVEVVy/WsYKQHEI7Y1SfF+1T63YJ6i6xLNUoWywIe92EFnNG6VB4UnLwqcs2Yke
7eeuNH8YioB9/nsFOj6RxJOkJoH1MfhNrtBLWWYCur3fJH99z9kyYs/ebu2IDMRp
Vbf1iGKZQCSpfw3XKepgoJZPIPEDGylpuTQ1GCwXEG7sx2ian/0zC38ZQt7MtrsT
IvL6P23+x0Qo9kIU44SOTH0WkafIF3+DZdbAwhp2IheAqpp/oSqc7+MThIOODJGO
7qabFZ0vC1wn2yI/IVNtEiFKX/dSZq8wFXRMSwrsQOOoy6D9fqOm8qywTQ85jpun
XAJmwBejZZ/5dmuWDW5lKrCqYN0fkLHrOKj1Pe1Jmh1+NWpcusF3evIv7/kmescg
BqBm3wzDjYhDKLhBQmyxdkvcNfcA28CliFDhJ8/LMvG9OUkFWyNa2+q/BFl4u//B
wKUGV8PTm5GgO9IMqOqEMDpSzsLlFkoz0dDlI6323htBPzRIKLMgWh94aItkybQr
99k//R20Wvccf40VCyW3gF2gK/wNzGTXOJPJnGhyG5DH8MxFpvfdXnUzmT2vyFUZ
IFkPUBUKSBi91syvkHkHdM0WSW+JX/0Cld1i3fFmnKx/kcVRXNzM+lR7UiBI8xZV
HYbEpZPwv7PAwTHGCjOalj2RgrmkQl86N7ovgPQshx2i7m2z5Ze4BWV5iEA9NZ6f
pXclyUIf03DbINvv9Ijs2LVAvlIv0E8BXs7tmWRrK0tL0B1RfiZb/aua5Jrkf1K4
XNdqHg4ZMSgF/J83UH0ILp8j+9Sej1ue2zwnmwSE01g6C8AZ/2sjQX8aU3wY63MZ
Vs6xppNNU//5svSv5ehthg7JMhmKbkp/yn6MEQ2hhvqMAEd5+dK+fCwm3/LDHdsK
G8zig4SMVK9gf3elRXGYyRAmrd1BipKUQErRIGjq3vaXRAfwqwBn3Z1q2sv37pUK
DZWYm+NH6w8dmAz03DM2gy75/TK2uTMkcU5QiH9YdBcfH1uQBOqnGUOaJPxmel4b
YEAQnlWOJ5uQtryLZcfuUyaOnWOeVTkIcCfF/nkQz/XmvNm8ZR0+ZB0cAD6mGySu
0RwO4u+T7CISs2aXhn0VivyDFRRc9SoUWSTySy/QeMq8ZhV32bQB3GoU7Uargiec
jLre5CaSW0gTRiVO+p6WaUzBIUOQFMVJZ0w48h1gmCz085qU+5lZ9dQGqWekDJES
Cr8NzIM8L4Nr2lAhomaIG4gDG3FcJhgDfXx6FlkTLyl51wQNdwI1ecV30UyLXVCO
W76HaET9WhqfjAHIBBbPETyzMM02cHGpEI2vwKpVbvG4yKhkTbcGjZf6/aS4k6k/
7H1Sx3pvxTNCZhJK/oHrZ8tVntHNwMwzzu9mpbRCSMqzxaAE1PHl4kRTXW8Y7Iru
`pragma protect end_protected
