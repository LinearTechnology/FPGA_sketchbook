// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N9nV4BV488mz7vCRndEwpGZJD/YZFyyXMTjL47kvpkcSIjjeC2LjWsLdsaAaeMgo
f5tiTo6rs+HbPvcUF7FWomQIVkbiNXtuJfMz3AW5/ihm+x5A1s42wzAYZI100saY
NsGoeIq0MnFvHtjyM4t0YwpO6JXDb8BVYnrp6h0rQ8U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7072)
+3G616YkNrGiq6juOCGPnrzBrG7Zt0Cs3W9IpSjXgiYblGn32WPwIfQyhBoyEbR+
r3tz+Mm9Ilm6/FxjEiH+7f4aEl4mviv1QtY/XSUIHN6wnk+L7RRN/sANlghCkuye
YKaDQCUEzuA1bjuqc0IpLXPIi5LnaTD0KRqKteTNYuEV5dharupcr94Ycd6QwzNS
E1vGyNohYWVgOE8sQvD3NPDIG9aN9RKrlY/P6SxxAahA9+RqC99biLheRjRf/uYg
7p4oGaIxiRIphMwnFAhFgUXYg+6l41PReaDYu7tF1ieUiX4Jlo/ow/rxygz1IVpf
o3CtpKvuxuJ4DzOYsT/6zhMeyAyFDxfxC8EkExs6lhJA2Ws0nyMw2LBZHHg7R51f
P8qeWCSVI1b0fBKfeX0BkuIT4CG2xYuUehiqYUeVGEcH/CoV1VEbcbJ0V17HrxUd
4z9stmqL1w/uaPK9mTnpg3F3pRAySc7O9V4wSQFrfKHl6BsOlyO+rUYMQSa+7d24
4kjmFB08j0bIoKWPhAlEZ89acKM9/E7O7gocrveH5K0Dl2JMnQuMF6aUSpFPSuvs
ZBy9ig0kZNFUVcSUFosA6UH6vvl4N6fG//+SZnqS/FBBsSzuiNlLrWGWVPeRm+WK
khuURKo6ytd1K7sTRxn7/L+6Rewe3s1PDarSfdMUJY7WtRERhhcSGFSJShva6eHQ
VGw0lBpobo7Wl9VhIa1pdlPcbWidZB9FipBODT3/uKnYDQlalhhTtkEBCTqBHMf0
hT/Fa7oi8Y3ldsCggB6+iA9HAXvoQpzkto4WTLfgPFuHPlRSifsKFeHAeahg8bvv
vm/Fyy/IeEtMT7L6k68c4LDCDp5wTFbY7JQrGbIkr45nA7QOUyl1Ql/p1aWJ+e7L
cObHWKrpUVRJqAk+0W+BvW2z9mh6nNgxg7gksjVxgovMtfgqoqSZGuLaqLzKsekR
JEH0+HGnuYpKbNrJAc3HaAPZ9tPZ+jHX2snckHmOB3rfrIGJ7jz7oSFn1jqLQ9n+
vQBpCLKQTiOj0/97xe8lxqGwQLOcnjItnOIKh9pihqL9qSoSetD6yDlYN9Ju2zSx
yy7CTnuUQHjF7LXHvOm4FUs140On5F2Q63kklzFqYzj/1mgmYH+i77j0+znDQCuL
0CqtYPa5IpOQmaVkQ/Uegv4dntQa6BOiTLVk7F1bghQJJ0t+ahyNm6f08KCIZPI4
gr+OAWPtO2wloCmXZCIhIB6ThMBu1vU69cwB7GxLf+Zeyjm+BvwftpC8RiLWENUL
wVvDB2qmJhf6E1W6mvv7PqXTRQEebq+1seZPNsCbubX+BVshfjiEwymfqb7Xke8G
CUxyggivvsXkURBzFzjf8QwzxeXhq7wJHKvN3LnBEqYh9CQxLa6OtnpxmGPjeLcO
/VdPdyjjYqlcmOV8I0U93cnNq9xOoN5WA+V3j/ZDX09OAfR4hZI7A8vg78JTs+Kn
FBG+GXuiYYiZntE9nprZ4rJRbAifo1wbUR+rZUIfAxgCmIZQ9QK+q+xmMNMztIbf
H19QrGUTrFUkFH74EwDUY6uzG41HntORgtYAujZ6y0P8dwZ/BStG0ZRhtQA9eyEn
HaQ0bm9x2Yd9Y7qAWiSs2Lc24pro1WvGM5IuS644/h6sGE5eBNIKdegPwcdaCf9g
6qO0TlStHcBU17V+8hu0aqN1l+B4woN6eCbOPTJ533MLD2Nkwip+Rzh3kk9GMR5l
TNYiD9lp6gFN/QIi6dxslPqqxdJPcxQu6UxbZfL3BY4Sa0GCmippqyE3wITDbw6Q
xu7q1UPrJkhEc9dAPDZZwNt9nREhoJr7FDra13AVCDzaklZtXfsvBbMZfUpJMTPW
SaoRH3o17PuPqw2EvIi6n6CGwE/yVYi8SIASbkReF2lPTiEkzs/KotHqgQcvSB0g
e9R8w3dNPofBNq7ZioWSqWH8w8zJlyUKiuoJBhR4wLbIq9yh6VCV6iB2Sh8BZTK7
aaDN83NJxG5sT2PTuFIH6gRZ/r9cxxfiJ1Rbc4Y4J4VhsJKgKWen15dsLPyXX3WS
jCjEOYyxw4ILF+tYG3uMBdW+jIUB5WjK3LLBE04RG8Tu6xtN2jBXv13tWc+von1f
SygG3ALxfhAqyPX0ZG2npi048GGYmFwa5rr7Y4KLQnSb4czaZCNkpKQ6MGHgq0g+
2xR+nYv5ypVou06p16Z+vYXEsJe7ehaa2mEvNp0umdyt73lLXYmET0suqyDN3eTa
JGTzhrh60+lRfQ9UGYXpmaXigXQZyYvZ6RwoLXzjGsBlhZ6I5OX39tTDQeqXzHsl
LSloUC4txi+AoZ+6yRfxIMdcUUySF2OjVNmyFt+8jRqx5ZAcjyEBUQSbwUrnA6JU
H4vyXZhvEYck1YxN+/ezP9TsQM5E6s+mUTFBkIqcxFu6JIcAqUtV6sXA1dCbkBir
aY384hiA45sbSFp/GORQQPEkp20/cQCIX6e7F63vxCLGD/RGqQkimp0f04GTLUlw
S/fL1xVbGrVaYW/bKFl7pI1N8sX2Axt3cI9v9aotQ15CebQsSmtoo6j02ysV41gc
seoLuTXvGpBEKLCbrVdcHvRT/l6qDeF3pNqP/fvop9YdOTa8P+OsX4I7trFNJXzs
rQrlI4TDmB+fluNX3igG+i764VCDgOc7HJm4ug7pIQ66WYBKpWUQ8RTMXo5BGnOz
BSWQ8KoijrNhWiampwtOJu+sKcrzlGrvY0NlcuZAEDm2ADlPFOYuPstp/rHt86iL
zs3krZ9emAvFIbgDOhk5eMq2i10qtBU184jIvUgKisWTCnRSUUXw2UQXZ7kIAb2k
+LPw4akjsjFoOLONC/ezOUuilRYTtjAI5YPlsrbAwEahpTNT028yoxGCEGFJ2bMY
BR3bC1BZ4WT8284mp94r/xN+8z/WjSLZiQ38Du9XFfqvwxx2YmUKsL/X+t/n7apY
4dcE3/nHw/887M38rV9PMk67y/OOgqDQPS6lfrOz0sKPXsCYzPadRrddsijFmH5Y
sCePYoMxi6I+AG2H7YQnEkjmaFetmhLz6Mfxh9oCwYV1QPRmlh5y/hmfRx5FSO+L
NPr0Me3/yAK/8xg2hIRJ1QV9ecGA1ZeVThsKN3HbdnGN3dgCfONb98aqhco92Jsb
GZyGs593UguHLZ/rHktd4n1qMqlEQnXlNe1UboVVmCdJ2qXuIdD3wAWN6qOfEHZ9
s5J2jUmqyMYhrCtayUtmytzAmKjh9ldtPUte0JuNhgLINC8NvZHK/ko6NmrTImdG
9Szc9Q1D5msSxpyZt5xW2hBM0HeRnfALwJESIHuX0Uyl6LSw1wof3aRwPxP3LcIj
T9n2ctBvsbPjudITmDwewF7GiXBxRgTEAYcs6sWgZ0ZhZCNhZN1WZ/PZzcQ6TY0F
egKMDC370mSUkjXA6TB2uE7TZ879wEAzHt2IzuYqYaA96I1NuYmRSm/s/rCopOs1
01rY6JGTIvGJlcnRiF3CXpmqdfOU8jT31PSJESPxwUswb9XLG/eimGN/giuMro37
NBkMUCAmxv1MHN7mnf97KjKhW3glGJSK3aNF8V8Jqv5xTt1ZARdo2YhXQWe6TU7i
pTAxSxP6Lah2SPNoRs2YjmoEm7RwRU7xHEXniYXWPxTJEWzaQTkRISEA+U2oDMoK
/EdKDjR7DxuMyMz3qsHTuklnCVaKCo5UMA8dGmmOdxXbMl5HpvHtG1uD9csKsDXf
88S8P8INnpgFaIg21Ypitv/wu/9dmxjPyA7G+JR6BKsDvy+trfK/t1IePLlQE+h9
bV5FsfiHTTHLUiB+FYNR4uZ6JJTq6y62Ihc8eJjIlDAO2Dg6k6+fQ8jplQAxMdjQ
j6ito35vYhIK2Bw+JdpoPNzjO4wjFQqCRW7fJM/QmFeiIBiIcwm98NEY0iErsG4N
VQ/gnWYjmSV5lID15eNskx1dXrcXKMFwAYTMckGoIY+iQb5AZd9Pk+FZeAeIhTmR
l7y2r2rfL8rn7WPCGZE8bFCe0Qq+mnTTMtxu67c2HNEsrFT+yKZs/s78gJN2YuPm
pD7gLanRelcP7wRDF21L9d5daVfH9FkPbopjkpteBWqKCj/3IsRJncTmKj0+e4cS
8ROF1NEZOKd5cUL/jjGz+3saEE2cND1cmXENnTsnRoR9iD/UPM3Tkov919tSqlMU
/lXa8FTX6cyZJ5uEsywWFpd9l0XYbo3PopHpXajq43TuBpEx3fkLXDmNavvsuSuE
7lOohhk1VTn2qwlAw4I1gGQcoUFz7s5zuD7hrKcHkQAqPfdocOJxzENOPEvI3+yr
BPDCOUIWFvzUJJihVhjioNNaaNXMnxeWk/sSFt/UeKhUctBeSCxQIMv6mWAldqJ0
JiIVQDMcXm/voUfTG+MFkksNgcC7vWKs51KKHEEJCLySnx6tvnpVuMpTL5Q08oTV
QdAatauadfPwScqqfuXoyPb1cTyGD++XcvzbwKNkGXz4rvK1HdmCWEVGQDYmZYNL
jQ/cvNVR9AVJdV2b8+jEpqtqTK5fg0lM8jXVcl2FoReKQwxlwLmSqY4J+6DAz5AC
AWVzy+1zuA7NJcY1IPqmN7S25psLmWaCwDNAMfz6MOwqPkSJTpA+KgIW9Vc6oAhI
F5K3dhLxmJs7DsPpvMfJglwdehaDRMflnKUvmtSfLxT4pH4O7P+/Ev0zbS6qK4Uq
zUhHdeV3CREgxE/CR/NYr+HEVOI3sFhptxuFqOhQsQGu3v/BhfIu1/HSQI1JDeM2
rQVNknXMDd5yEp6W/4T6Be8ojdiqbnciziUQq1FK60lLGWY8JwNRXV1DMdSofwX9
6St26Uybb2VI/Oe/wEvA++SczYDztG70VLiX9TaaeWs0biEDg6boGiAc13Q2TBVK
1Tno4oeLIcBLgEBIIjMcLWzozabCGyv2k9qUYQfPHOPr6WwyspIKZRoNkRoy1qA/
EMWt0acr5U3GpwyyJsiGSdLefZth5erwahv4uncq/zPFS8VN8EDoNGVwXqmENUVN
7I7Krtvqru9ez9y85RRd8k9dVqOaBldAVrMGMcKm3wFyD/oVHR3KCLVoDkgoZ14u
PIV4NTMfxUumkT0zaxTDFPZbrih4dt8O1owFDHf00KIUpLPPTKQIXUqp04GRFUBB
HoHIVMiQJ4sSMkqZmsibwu5QoHADDyt+eFFpiNkwiK40/ULNaU9H9VA70RM3CNpv
379BlEzPc0T/Zkx72W03Z/gqo/DCCr1rfhkbvXF2kRG4d8qmBDSb9AddE1K9wIud
YW73hohOioGj6ba0jtMAKDBnxrKVALrOkqEjIp5cEKCC9IkvoIbPBAzxTt6EVpst
ZmqTmjXNf1Uvpnmq/ro+ZTefWixxqUg5XxBPLO1VPHHbe9nGM+UoNTG7xSj1El8h
3DGDokG/N+k4KKTjOJz36ojJJF3H3D8bE9GTdwvqgcPsktl1yOJj/7jGquxLAQH6
3NRwHIdTE8t2xRp7NgG5YRAUVyxibamLOaw0TR37J9nDPASl2yE+ZUKUdyRaMcw4
Gy4iSKwI0CJtVlYiozKgxaN+2P9ukpUT/SI+I2ch1YCiM7C1RgJQ6apWnjwDoNv8
BsSfut6qW1fGeBiCEhgGjpS0F4muSQDwJB0ott5CXrHazaYuheS688wLp4PnGZZ2
sS7QH+qraPazzpHP6EsfEwTMoj8lOdD2PY1myIp2BNvc4FBpy8MHR7z69nDW4Yei
QgDY27QtBZtLckftnJsSkFVCNfwNBha3FdPzXpzZEX3rvNvSGQ9Y2V+dJlQAa3Fv
QEtKNn+jo1EbRRdhvu8KaUKdqskwtRg7VWcgqWecGy6haZ6Xn38weDfMHZgsLa0N
ONtX4IUQVRY1vPDzzY7pljd0mUVFnk/x0bzN4kdo5SNxOzMNidzfC/ThRoJ+ynrM
5QUYqOrxWxvP0RQBWmfc+kZdTqqtDcmYuubH/c9LwXaGdt8boMKeImSvobRs+1LE
Z1CXHQ/M6J9FqfxyIGvCb8LpJ/mBYqlYQIo5JVICiQdLyO/bZ9INx2uc7+wFvhiR
/l/Vu1FC8GPsoNbXaDQVfVadOMhKtbuEI6dXSO1rnxKAKWxjjwYIdP17ZLhoXZZf
aFPYHc3kU5VhU5oLCwEbEbEIRke4pG7NXAkOHFsHfrQtKuZ9rz9vp6DvPyQX/BOk
11h8FOZbOzbEbrGX2xVPuzyLifi0IkVKs+fqaJlq93wdHKBhYNAARtSDtHFUqNEQ
Qaxj6C3JhglRQpnDe4bYkhfM0704ZFjgofSuoEwaEpWPbhPGSFFIIrHckNkIXYR9
vzp8m0DOgfgehzrfYoo5t0R27ch41YIPQrUClZgFudu3icLT4Iu22KcULYEt7zj0
LeN09/QVOtCNcXza70jyCeaGieCO5ntYYhssU8v/g4ZYpAP3PAIKCDvact3jcZl7
4t9epZwXFPvGRrBEKLyOWS9+5S1ALDWjZ0PDKPTZlZuSDWB6TOvvymGMB53NFXQq
B3bphlGKJ018JvAUgd28VsCOL1qhQs9d2CVA24eTwGZE8gZKmZPqdF5HYhCu3fG4
iBEfJdnK9rylAWP3uNGYkrXPckkTs6E+BDmW4HeFkRtUwVp5w2u2zt54wM1l07ia
xKwunTtcrdL4GojmR7RkRtz/T9ML7BypwAL8MZqqCPwREoumurmLb9d/lByWK8u7
uLaM+wTmZ55OCCLDEP0uUbX+26OhTCTjxNAGsUPLK0OdKCOoo5D8PQcVN98rA5wF
NIQHtU/8xq8HRBNcLJvRjNeJcJat5QpA0Vjn1RuKesYf/3asxUO20kzNq2dsM0wN
l3vjJuhFj7yAeAJnO+YYRihsYK0mScIaFuVKJxd+iMdD2doFYKEWm/uAkk0AbH7t
fG+bNQRymX3SmuPaXQoO1KH4cynougV1GqIBexPIU0Z/0q9xB7OF8bz9++DExuOU
e0lUIGHyjld9ngjrzZadVyVZYZp9LDwP1THWn6eTVHQ+SzNnb7mGTjZ5R1TbKv4F
i96nW20toIjLBfjNUGgsCO038qjO322+eXlUurhgJgroKIyh5nXLj2PcJGvxemYO
EURocWZOCQHMzoBtaeX3rQeMxc/or1NzzoMYBukMCJB5TBBQ3XsZvjx0EligNBue
+Wxl12mz0avkHkMTorN0/BSRtuWxI6zpDNoivCR9tAx/7VwM1iPiMZqla2RCPVsc
tB0h1y1u1dgig9qighsyQ17nDVtV+rhE4MLPHiuQZKIHhPLU4scM6fNf3HJwEq1r
2bAi7u+CbREXStar27WHdYqHOvzxoV/rhXecFCD8LlXTPGOO9zUebC1pEDzDU0kk
X1MkAw49j0zBxZsqqJqKPJIxnjBoyosLAUuDYPCEzlKbLQawX8w/jjkDd6dDsaza
ozFLH7Rj8wq2ijdpHsX5d8BNdDhCzrhT1C1bme3QG8ceZPyQUD3JOd0dL2+ggvTD
olInRGfBFmrMYtnqfJMwhKoqJrr1UYTqlxLF8STMSgLLRbHTpEkDccxv6Fh9sxg0
0RwUDui5wUb/wVk5+R7hQ36FkhXfUVuz/4v+qCoAkwk/ZCPvZbe6clAUFxBp62ZW
gjqd1xPdS5gN3a2SqhCLqelXZUWk0DsHz/+Wv4y60+lk2P/z54nPN6A2/vTU7Mdy
1oYvXSse6kxef+vKVKFBmIk2/5eC05qHH0tYq83lRf/8f/GC8KNehV+J0u27G2o4
G7THqadQoTZ/7emfOKqRuwfUgF8gDlE5Ioj/8TamGHGsQueHkEJobhGxv9dVar2Q
04OkZbkT5c+jCbgiTHyZ1Ui+C6MmAeyfejsKZV9RAdbkc2REIkgbGBSGcjL/5YYR
6VPppnWuW6psDwrBE5OB75ggeo+3XblCvrhb3QbBW5i0GYhs/y8MyjwU4BJTI8bq
F8tG8CmWKkIlbpGvB/dbq7YeDcG/MVpghWVTwG5I/jSyDwn8Hkg+Ju8jIiY8b8n6
DoLtrXvXJD3+6Se6d++Ca7HZrrZwomH5bL3YEvULueRxE0cvjQoe1DJZ5/GhLQNO
GNw2GjwFm5SBB4CIrNP7SB/LhSkRvVYWpmTkKC19ZtuW3FcNrW6aKACfxTMn7GgK
AH7moHVErEs7RCsSCJDl/iY5RdFVvlro0Lu723lboz2EOjjqJD1gmgoHZPLCE85w
cDzNVAiEtWCeVA/ZUM7urqJGad6EQDnP2ZssqiNU4HlmTnzsxucmF7gMq0SgNf13
+CvnPg5UpKUUWCSw/bNLG6LubcLwYTKGCWy9ZAOcUtrAYoapCEPpObvFwbY+yn20
kkNdM+ZrwB8WzqmzeJEG8iVFwzC7OrXwAUtZJpfe7ZZRp5IULZHLhrlXXtSkhvvt
TrNVXJpF2qEuE1xfF5dX+1vov7ZG1oHii1188DdvY44/k4l8FLu9atOk4DyA/y2H
R11TP3u61oGsv0VVD6tTcRHiamcJxF59EczveVnp37NKFgYgMjgGZcrgm+dx/OVS
AfpQaGxq64ocQ4kBJQ97H0CRiwSjXBIsmhtIfMqP+2b9cSPhUFN+LuBLgCN5fRUR
2xaaq+ibc1Lk/E4d5ofBtWgTaSkoSt89Bd04jxYkljTVE5GNAg3942Tk9uTRQC/T
r14VjWX08gTypmcNUNsrsg5bGbayEV6PvgErMQnPH0z7do4OA9au5cOuZOQvHDBR
+p0JZcb+dC2nKEiucxhGC53EB6MlqF7cugKnH3xGvQe6nOd2Dsldy95opQAKWEvp
tixIqGBT3p0te2T3BXUvono8w+XkxZtCcHEe1UYNnlBTqLjP+6RA88Q085FQAHl6
vXlFvGd2n6pxV7kj+Ju0/69RmCgoeRLH0s+EfExGm7bjsTU2mf95NuJcJrDclryy
pK0dDbepfCoM7Rlh2uQ2bxLM9Y+g1pHtkkB3vIyiiI0O7Dk0H3WhJCDjW1+e7vJN
fQUWu4ZkmyAsWqitehd6rDI2ZfTegswMPJNh34qIiT6FtSsHKW0kSNC0aZFu1G0X
sqZ9nGxAoB1FPpxzeXuMIkK3eEXHQ6AhDVwkr/MyetNuYKyW+zSTbI3iSn8Cnczy
GhEB3jIPqNhELuaqCF6E2/1tAI/7fX/+O5mCp77O1bHjIUWYAI6YE2RuGScf0iCT
B3qdDbrTcCCtrFAgptebMQbLUSPbL4XetsTJaoK+5DVGFJ5h4sQSzpWAXplQBnqG
N2OBm/7s8mtk2c7KyCb1RA4u/7dAxvCOPZnR4+da39buRQAYL3l8+Fcbq3VzOLCO
Z0n5+iBr+2ATCwprRs61D8hj5CgC8hfX3QrWVwby6Z2lGqBEPmgPpmQ57RzRpxwN
VWVwdbZcNN3MXAG2n3DLo1IiDbrVbl2gcA+Fp5ZGTdo4iDsav7gCKAgHKa6Fp623
eBsIDfmgB04hXkjBCWvjIGBBpvIeK+b9V9cQX0g+rggOztoVDwk8GTdGsCk13ECy
e+OXxdSjGhbphLHLX6sqWQ==
`pragma protect end_protected
