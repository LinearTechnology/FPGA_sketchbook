// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KIcJ5eJk71vNDYY6RMhMPcoy8jnRGSN/g4qLSH0ltYgUG9mgj8u2yUJRR0slW5RG
WjdT+EWLqC9OCdoAI14cRYzxq9dO0ytHmkZjsDK2ozex/rKGvTfQE9zTYwjyrzz5
DUb5NGG2IVxy3H/B7aPDMtIvFPSRH0PIvzUABaftiTI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5760)
xlBhzTK3HkNA32hwqqm+rNeDq1wPbOmOOWLEJFfCNP+yoU3EsBbDaRj9ew9pf+nv
rhcjg5lAXvz9AzY9zbh39G/FhvGJNYJWHz5VdA9sPcUrHArMMBQNPRJWRJLMm46Q
nFw2Rt+10sWKVNiywgxndFU0uJzdGcQ+gn8iHPFUKpIYD8sRDYpACkwNiYptc09J
wz3bO0w+fp0SWBiCtXHPFH4gtKip6NMLdo8KcX4tgNcqAeO2gJIZ2E/KspLTEug7
NqLT9ryG8xEijU2xyljBU9JV2FoyW+PQPxxyzNF6jRYGB1xyPBwGbZf+FeScYmWR
lkV+PliiL0morYCvSmnhauPv/0FLHCK2TU01dawBzFS/vbjCOPvTm41SPwFJQNbe
DURY1aYjFNpi/Plzjf3zYDm8kUrBss8SNZeIEiP8cmAsygIlIie40jpBV99jWUDs
E1p9BtOv2UJmBmx7XNQOXfYNp/n8tuP5uCJgCVRXyoSDIlEEC/ax+xgFG9MleaML
PGXaWOrkCe9w9KyIMYmQrvkEWDpfplbaQQ0l+LxjLkg5Hd6p/eHvcXIbWN6ousli
NwTgyREbMyGBT+cTEcwFBLIbUFBwTB6ZnqYWADh0CY8vrs18u1P4SP/w1dsqdDT+
gC8V0SgICuPNyCOpXN5iRUw10lNV6X0T06GCU+EoJXaYMGm2T4YNb0eQ8NHN+dvK
okrrpMtBj9Y3wjGb4oE6RLwYKGZ3gU70CsFwqR17Flt2EKclExpepm4VWk0S6Yb5
+pGJg+navcyL8sZMJXJ6wBF4lu0kEY9lZfTj6S9xRqOf7ls8sjtkcKy09MuC8Bxq
vmzBvZG6G8Qp5UKBwxVWCkCJL0hqidDhvNjKrte5XpRwOC3FyeMxYq3cyCwGVFEk
RJeMmGd0LsOwNKtCG/hWNQr6ktnKOiMRFHJY5FQtiBcPXVMfryvHZWLTOm7VlCi1
dsHij+tvFjGEd3dPyV/djMw6DycG1hrHyB9QUU88JQcFTPdm7dquc+CtJxkW1glw
nNaRIjlVwT1HLn1HKUv2GSRiiGwmHNsbS9i6UqtRxBw99VlydFxZUYTeveREfdvD
WiNZVMOwOqDrzWj0tA0du99ZCTxfd0807vkf9jVkK9wk7JfW2uCch3iUcz/foOAn
GFzA8G9z/zy696YlDC9vqHeiOduRsUOZxB1ZkWadyWbBy9G5NmFVULh7QKmpsx9k
ykL6/JClwiK9h/7eNuA/06lhjNwpHRUcszf0Av27ghuYhmCljkIVO+hDNNw8wT29
nX2dhkdDj+E0wHRfnm2b+DBVWfsyE34EIg7OH84syruoZQssVR5qPqvMgBXFpfC2
FkUVbH7bdG/D2KSj+SgeMZSYU/lJvP0GTxmXDAKuY3uEzB4FUWkXrUwV7fbBrsHd
E3rsoh8+Q8ijaPo+iebpdSyJOrQdY03dIViO+G3Xif6UtHa/4ENeNJn+01oJmrrk
ZG+nP8Tr/bOkF8SpLSLhikdlP9tBqXONCboeapYpG43xfWqOvoOTg2FHjsB88x7e
eeWuLutswjM7m3R2bBkbKx5E1Bnh66Bo8HDnwJXBbWbgQiN5zyZHe6VYbK0RfDxZ
k5/tU/Qxq/qNuWND9IqrJGGPPecNXP54y7/ck9+8w9C1AXlpwGYm2Ys51epnx/i2
K6Zf709+8r3AgqDEqUW45JIoOAMxhS5/QdUxpB4qF+Oa6CBBH0URVZrrvdJbOnaA
4jsubuoxarOCcj9UjoDPgwlKf+q9lYEjKZt9GdhijKXf23RkYHgaGsHU0xJLsy//
N2MqJWtMDaaoB4Hqjd2zY9ZTRlO0Lu2YSi4RFu2CGttN9ZRbXJn8wzaPLa5gdEIx
2GgqRXhvU9TzM1hWHs/FS9vjxL8bFBQ7jNYiJAx4RfVBIuL61IJJ2bpdxqAzS15t
bzc9xA7M60dW1x3Gc8uT5yWlZrkO6wEjZMV5QyChNLdW6pKcWTs+p4aQpwPynRPJ
3r6nKwiv+W1FrrTc9J6UahG02o7XYEANYyz5kisKzmjwMtpux/cXJlMQjljjjgL9
/szKOE07b3VKzkX2DyGRV4c70ExhElk+0+or4yxQ8HgQP74OaMnHXaQN4zsfHpHh
W+/OXl1MNuQaUfVO6D7hQbEsthXfIWZ0HZZlF1M4xQ5gZxfswSYfu/DBQvhOPKDR
vz1qcwx4h8+KWFhlEEEQPtpmv/PuDUwir5aoL9KecxPcAAGQBWz7Yq8qAmVcjWvC
ZM9173pDQbkx5052YwQxWfwQLIHxjM0Bz1xkL50YESNg38ncp5snbmuAZzofxbsD
a+X2Qek24sssaxm7md6Ov07JgRZPkDNnIGuXb3GV25q2kmeJHWFu2JrNIcooaDVb
qSJdrktmrqiue3hl3ODKGuHk3eFp3licIqtcNXW8DEdVirVKggCxJPcfWrv9brNT
/9Pc3S2Iayf9nscy1EyiGLzrojBlWpVMweKyPVmHakGgpE0u8KSW60KUC0pChf4Q
BkngcEHGXT84OgjnpwxGTLUzqrIhllG+R4JtTAoy26tdheyBTCToYJF8krx5BGfS
FDha9IIk2oUT8G3kLmMPxdKJaxBWveiJZwo3KpHtJReK2D+E/bCL9LAXOhUk+Aub
6dTslDOotPpnAXiYA+5QhBNaPHQxbbVOzaww/OHUa/Rs3M/r/d1rUvqOm/oAWgA9
krh+pNhIx/a3pYDLh4RN4NXsLPnEowLxzaaOUTY6e8oQHsWXOYyJHsWImveIqfxi
oBV36i/xueWmRNPFBbGmVJ3rOdn8UZzkioMi7J1z1egT4j4+vaAyk0R4zSysqVPZ
l+12VHiZLjXPdawklgmSiuwP/nDypA6JsIMwjY11sp1tbsDTkFJMmxpmsrmmrdY0
Ngdp152jRbnuzZaa9SebBuzF6YOS1lDK0uDV355eBKd3u3ay+lE7KuZMRCF0jkLm
hWUr2PRxvpmDwLtRgc3zXr5gx12ILTRPtTC79LQWSZhjuOR1BSZoifH+PggHhllc
DhfoWAFFDrRgQZuPz4yuVsHh1A3GhBRGBdACX4aK/2PR9jEGxUQmzWQVoFrpeK4q
t4L+RcE2WuWT7pjsr/G0TzGXVcSja68O5/yCxGUmmcVn5JhGiZHV1nbPzhREsNtN
kHGoCg6/FczFgoLnj07Y688vuTnw4fCRSLk8l7oWc84K59ysscZXtUgrMCSmdZCx
/A6WxmfM9XzczQx0KuE3eDUp3rPH3AfZj8/36x9T8d6GKGmEmxR50MYWgm3hiRx+
1+1MWXDqBa7ze9rgAmLklIUXbD2upqZIJpco4xCHWFdgDuwcCjUH20O2vriZJXCp
m8e16bPIZM9Kx2CcotWFZWEUH8kMk6LaYkLvgXjPbfqKKmvUJG5Q0uiXNPdX7ZgS
w5fKHet8SEAd8JKk2jwYnePKGfDOwNIAgvX4tIeOH3zRAic8QbeCL9ux5wAKu6Xl
XBWp7O7hg++5k56qEznjfoONZzsWwjTQx6h71nsmmimo/PammuAefbKOOn12ml9V
xh8grmdQhyQ2oMbUem1ifWbZtF58Bx5j0XcbzkDAf6ANZY8MQeOlwvCgmbF0d6KM
VYvyYF6IpCfkSJUMWk9tgH9q8qI0Mieac76X/09ugetLkHjT9AvJFJA1za4NL42N
u/rFvje57MQ6CEpa2ducukHqrl/4Y/3UExCkD82e+/XvPHiWz50IIsn9sudbPa3+
tuQTd5pzW5RhDSIKoOlFkPxOHrPEbDRnf9xX9BjHnq93zFwfeP87skAovzktzb9x
qndQmAMTakv6SJ4LB5RzJQBpxIdpTYiSiG/iRJuvVYcNK5wDkFEQoCiFgudn30+z
qOT5wrwKBJhX6l/V7GzhO7POtfY93K8FkLFVpfXx/V7zELD3FXm06EdWsbyLyW+0
1/nDx1QfUERQvNn+KBqp5VUhRrplzs0CqLpdf1no9/sXZjFJg+Br0Xv2GMn79Biz
Z5ALK1zz2wzjC+eTmgqKweo8i9LZ1AQWMf00bj95URbjUxvnjkz1XiCNxOUANyk3
11dK/b0pZBrwPamdNkhNmmZ3BGnL9+SPXzVMlsZPBOWp6kEbwLHzaFm+RjXPHW/9
V5qseEOc3hYPF9QesXRnXfpnNQlDBpZy2q7zd9c7petyjbIlvSbBX9pV2KnPlexu
8bcOXd2mt62sUIkppNIdRL/m1KS/1s5w0ZCfGhRF09qA+RniePvooHrTw4NYT5JD
fAlMtmRi2yVUfZ+FFXCJtfvyMPf2rsq9u5Z1dgLFct+Gh+oTVWrMOyuWZWdfRZtq
4vsMIHzZshbmqNJ3Sk1G/22/k4gHhwP5QuRic2MO0X86DLp39QLCIApllspLcFMd
IPEkqfV7dedMoy+qp6tGLdBi1qUZbR7LDHmi7+55dx1qwkKzNBA9MR+RfTZOof+2
y5RmE2bmppV+6DzGqdOMo8u/h6XQdc7aI2RJX2ppeDGjbDAkRL2HUB3n5DccgiMs
rd2QfH2YBASOdZVqVAIAUmxC53HQrW8G8PR2JhLmsaFfd4O1wFg1pxZC61EgEURA
gdUyPDJH2qFdn9BpmCF8BEKif86kMzu7+pHZDKPoQHWKTyJeya4kz7kFNBsqD9FH
JCT29TbUtUafkLfiXJ8juECYfBLRkI9rHwqzNDoYR4tppKY4lNwtwvfV9hsCGDND
vc8P3zI0+YK82EHNymJiNYmr4LHEl2zx7K2fZVucg8g9bw6/AXSrJqh9r3usAmZZ
gdHQu9stGwWSCe+OIbokpvfPaGp7ED9GWEyMlXM8hubToNVCje3OVhQHoJPHMMvm
jfUu0nMcQ89Fq98kOEGI7D9EoHZ85zRnP4eoNGLWqetKVotfT8uGDJD4vCVdhgx7
HtxRRlZU6JrFLRXpHSUvrbt1YPQyhP0IN4M3SezZlkgsdeP+ohBb5vChD1S11Lxu
rTPNXRrE6Z1v1Ovb07rys9KJqXZ6Jk+WOoaYcHxAAP1tUpsNwMJy0vLerIE2RS7e
5HcGNgw9ytygW57BQD/OJ07rpi+U+kCnp8I0utejbF2qNnDyRrzTiJ3FUmeDUfcE
cnYV9zLVzAUfigXYEY1lGfzOZYOUShTG7P8UFAtQdpGF0uuAwdd1MJtcSpJKeNj+
aCQyTH6gr33FRbu7VGBLjtoa3Nl4GxqE2/lLE5FZ4A4Y1teKEMqUpnYxhGjx/VSX
dx5Ku5hYdeTf38NZ+Q4z93kX5qfnrbaOPEhMQKLqLWHecUGFFZPVlhywvSVZVLDR
COl6lfBlJEjYE2jeGg76vXmG3S8iFSwKIoofWWn+KpUHlRVHlnqi0QdtI2DAzZ/v
oukzOeRkVT3dVFfCF21XkEC9kkCFq3a8Ly12HnnPW7wNT7NKLvdL9xc2p3rQfvPU
Uva10+5YhdmKQTIRLGdsbhJnA2KS33LxL0tYtka1otPGaaGn0LTfVh+ddZ/cmd9h
Nw34Bkj17XCoSzoPmIKZqYj0a5vYIObbVzpuWVMtasZLby7RxjWe3XsybClK9fFF
gYLeWF+Lbm/uj9hcbK1QYpOPExKhgXeusMghTXOJf3YpLNN3Uvn5JePZTGIgHTfj
eU+mZQffc3O3mEtA4c9+ZZSYxQ1/P15EhMafLFICU3wTA7sdBpjTaBZyo/LGhBnK
WUTVeG3TS3xmp7rM9Cr5Aaaw8jpkX+NCSMyVLW39Yt4DT2gozB2R1w/UI9khiGAD
48lGUWuJHCXXLhxWDzbdc9vbfa/KP8Urktz+jdb+W4E93h99AcBZpy+KGaOsf/lh
uWMaJYIdF/vJi7eXDwZPwK4llIcKAqRbbDpoKBsQxwqTmcxLW22K8sIp7suW/mOH
pHPozgd9neC1ap23R0ivZCOvW4fLci1/Ey79M89HoBuL7P6e6+0hKwH67K4/9wKT
YBajhE26TjUxwtLzh6eJqV//2jV9wFZK1IwVf3VG+AImjpPUtkE1kG75n1bMO/JK
dsuFU7U/VfcHKhoCELJ/B6g5YhG+keK697vkhrDTpH5RSliE1JajNvvg+7/9VxWo
EHgLOj5WUQwcIT2JfNzblAYjjUe6CO0zCDTfGuMswsqJ9N8pMHtV/wvOQgA3zcyE
BXNX6G+KLZyo+dDJvdplCnK3FLmRcLPDyBYVsG7nYzYKrpnD94fJKO3YZ9/7FUJY
AkLWXHk4VeLIZ2sPOMLuG06WK3RTi6dE0hiQ2UeSU6CadRWba1np1NoFBv3aWAe0
IVX40x8RdF1B66rP61J86pJ+Q3+1I5z64cBKxQcLQ8M0HHi983LS23IjHpo0zWC+
V5nyzSc4OStlmiB9nqhbCdk6oD8YFkUtqIlXSmvgO0z7pNQ20M8SjQhZ7jnFVAnf
owlF3lpKAUWf0KFeoLPD8qTULMIfrwFtH/BM+LdXqvXfPQ1x1BIebb2pv+zsYHgI
afYxGp7kH4n8zhH5gGEXJGKZq0dgx2BKwVjbeoPNOdAyLswxcpoFeawB09XSJNRC
bSeOmQFyzIqphrVkR0LKCLvDUW7EB6EUP+Y4Ni49FgJaZx1lC1yh3SirsoAH72GU
hl+CL+HkxpSSNQub+W2ivXPSIB/ULCgMI/7cROO9CBsLKaAc5xVua+P/E99/veuG
jiD6NdGxRspuCuwwPTKEn38HWAnX9xeexXxCFOY9iSkGQV4tZ2jU63PvMX6yI5JC
kI1L6s6srjLEi3XPGjarSFXmuccrYKoCWSJrCCi6ZInL46NyadmHm8NNYXX6hUeb
ZqmLUhW9GdlCXIl6AGSjmXjWGUC+XGcDTIw2gLwQ9yn+NGKiVJho1qMGVi87ftMy
lIsCSmPcefHpySzFdCz1l2FoaTqOFYI7KJWaiRBbjL9RFEJ7W6MLkmEKD62e13Vq
Wux4EJDIY5DYgL/Km8wZ3Rx/ZxP40hTcnW02iqgGAtxga/9n2qeK8ewtZRPdsUAu
qHW3cBbfn5nE/QIUFZbsxFVgOaR7nKngDf3ZueTdr/ivDyKwlQQsiy4ObrKdlXEj
GmyVt/RhQM2lciJrcNVy/CB0Dn3n90dlLf1FMQ7lIxx1YHY6qHqIf+RawK/vVA01
IxCuW5n5tQ9aiEBAOWrWVdHrUvbzqVfSCtfsb7tYS5Tz7mQVwJsX2hj0aISByhdo
+Z4wNnUhlisQySZ20R54jgJjdtSvIOcXq5n3W3aWtXbt4j92M7sIOKIWHQkNuPDo
iBToc2XC+8u6tl4QOXdUT18JmESqoZ3aWne3Vb/y3AGV91CQDWCIG/xk0iItQ7Ti
b8W5fWj7GBDg0zM4QiM0L7wQWwlRGNuzm215+vmwkJuZer8j9sTngvf+pUHKlzLp
o9MCfXCQHAjJPBHKqXDqihARaJvi4N7hIN+ucgFWxIZEsZjj7GXtvFYttb93njYP
iY50pydQLKa4Z1MR3gUR0GnaThXJc3CquqAFrshRAH1Utdacm/VhbAH5siCdW33d
FEp894bSOno5EjDb4OVopyaKcI+ciA87yaMckKS9/I5tn4Z0unFh1Wgm8DqpbskH
akOwfYKzqhooMcMoi7bHo6Z9xwH7FgWWH+MPl6gdrxSksqG9GCCuPC4ZWiqimEwY
2basxJ9lApgQQV7ZJiWuOVHVKlDErjvg4Uo6e8XGzfpfX+qSt2XBTL/LVqd/dkRE
8jHBKdUPSODKh8bw+DTFpdlIQ3Mk1+6X9h04eG6siKRTcAueiwLq2xqGs1rva6A4
`pragma protect end_protected
