// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kcI1RVRmUqN12EGittcsu/rFYBHp7dTrk4aGXrEUKfMFVWb/iARMsRsygDhWdvri
F3YoJ2Z2CJRHT7dAP8AglmQbvlLG7ngIgBg+ootlFr9SVshU24ra2Azn+URDJrgm
P5BSMdRAVESSgxubXVjrEjRVm3uR7zFMfT0YwQIjxcM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27824)
IK2EPx/mySi3+PoXwGYm57K5Zccy7cvwWBo0g0/HCGYhRxi1wvqcqN8u02owc/bB
0ClarjHtHykFwl4vclU6MTMfMEua2rr7ewEme10tCwB5y/BrWaSH1UjCCQM0iBMc
rTFURZoy5b8kdoQ7JK4ZZ4J2HZpHEc9Uu96pBhWOheZoEd8D0HAI7qmsyaFzLbR1
QJlEs6+CT6XPTGDKA2lNwRBsZADUC7LTPlGaYdMYyZGWwVDE6Qmzo/gHbjYDdFWo
gosIGIrHjfJnzcbITUHI1e7QychSKW10oABF4by6L3ZYcUEAjXLXQNDRyqbSmELQ
kZIVSCvJu9Z/YAtmEOoTsWfiSy5sL5k/N/cSeClpYDX6M1to4upsAX3JB1l4OPNM
l5TwHNkk63oI7JMVAc/zRBQ0I5mD8foe59C7nFGIVcLpikNy0fdwU3VqBFYuTa7u
PPWjkMibVPKd14YKtjXUiUIoq+5UsxzJoe4xuUrtrkIG1851KOzA4BCvwKyftCxp
k5XKpd7OxRGrDINJ4iZuQvZXlWxHHZ7mFOlNwvfbJPZRLynoWTWbjLu5Zewm6ZRQ
wN4wnuhrHDgG5Y12w/qrhuE5+v8pSc8hagNSxIfwr2RfgB/dNke4oXbi0OEMBhSV
rHZTiKb12QkG4LtPqlRp+Hbcbv8AaIZMW8fqX23RS56erSQHSn6LM2P5hDcet2SW
e04M6L9/Y1W4+1IW088Z7nTLGF3HqANZGuCwsTYnYv739uJjC3zUds53mwRpSNQ4
+uO7KKCZN4Q3AGlWFmU5g4JTHgR4uBevmSf2Alqv6TTxlMmZnZQj9vLTRNQOWphI
YfWJuQBYrQe9A6D0eeWy8FW9RAJOMv/FFyeAcXdZDj9+n2Qn/fx5YCN5oGI07DKO
g+cPMy2NQ1RdP2XkAZS0V87RWaiw7MltAx5IyPvaFfOiwiVG3S4TU9APtX6nlq3d
joWpJ5ysZvdSdup9SMI/9ZhHRgsVFFAsyIkqNupBUrs6jJq8mti2yNPaGRaa6Nj1
GOVPOA7AgRMNtu3nCRvaPsRy/Di8FdURDe4i5srBiSNbTcHzN7OcA2vUoqbNFre2
eitFShXo+VVkkQyLvMsWAOn3m54XkVm3/SCyOkFq6HflwC2RGuMAlczN3CifRFm2
wjIefL8r2tjM2KRqL0R3jBePWGMaZvODGAhkuFsjUeNh95gs68JbM+W/ZUiO+Pxt
YToOLC1b8FZLYPckj5jwDnYNcUTOBFBnqqVeKqSOvfq7sKtc/dTnHOxaiHouoPZt
dyl3/x3dj0IJiT1CvfIeRBk8Wv+tPVYmnaQC3HvI5NN2aSzTEbTv8OO6NQ8xtKmq
4FqFd9fU56IQbOFFrDZfKgCoosB1kdQUSKBd8v0tQT/UHqa8YNBvgSkrCthOVYig
Lqz95VBkqMsFHH4/qXRRuVV1XTCCAt5fVpkSGFFHNPdH+bKs0nTOOsvdRpW4Y+p8
cV6d6X2NTGx3x/gFndwDXusH+W4ATMWATxhEY17QQl7iZVYJpfDMbwBMl2cBHPUe
rCzD7q4bBFKmVybEwLLYXupgZUjU3fCLx2tb4R5B5xsQr1j52Os4lclb812jSDI8
ZbqpuQ8z2AkCVR8xZ4uxub3h7jsh5Z4WqQW8CoR93CqoqgGsH3xI+FbKENFiYgqB
DamM7ewqMeMZbrbqHUGPEdEK3PN/QUFKvm7uq5hi7TvDL7gyXdx7GK6QGrIh82ks
Z3ySrpNFfW0KGsr4uBcrXx1lalM9d0HVmM2f5ka4VoUyaDkimT6Y0hFr1qasXsYZ
C4q6SOsFTkRcwDQW8vGSEw6iug+SOY47IICJ8kejgr9bUv53iiUMpuslWVyuRQI8
Tt3S5adFq9brp6wfsT/5MuaO1Iqw3DZMIjuwuJUpO9+GN3sU0zYDejudCyd7LIxb
0OhDZXy7Ul4ZhIpPlWvW8TMDQVf1hbhZKgFfMQWDq8GjF5s6girykgPqhz8ZGVCS
VzH16OLQ81z4crKTttN8TlG6AJoS20z+ryPWThoHkINvJlhI7FxxUfLnM+aoNkov
6v+eajo9FkUSNZzAKb8NsVvYkjko3/9/xhuhqEXvj7IehSdg/TgnHY4dcFXiPvKL
IetgnS2cXIj1kf7ThDIQ10PDDviF6Sqn26wZdkGFTtB1A8hYRQoNpzvxTnllKntn
a/5sLzD1y0IioX00d1JDKWerjabdpiJhohtyGzlvyRxeeB+snkQ5KaU/GZoaklsx
uSZAWt2OpN0elHAFXuSR5yCkOg/LZ2gUURexcHZAMItvac6odzSQaHWdUB5fbQY0
GDJmnhXv7GA5QbuMTkCNM3PLuVXRb56a9kW8TsHdxkOuhKAD/Rbj0ai9x3TY60J6
uWQ+mubEMl3592OZiTS0uZ+BZCm6JyWP2LmtvGhpVYbQyLOzD6fuDkiQgStNN7jS
KxNZySqo9NtmFDg7nhbUCM2TtBe5xeP/5R1lXCddJx9bMA31ZbC27GheMNffArW3
1LQFvfm4y+LsM9Rmq2qfohoLT0Wd030SlWs9e4lFmOCVwCTLLl0CZ1sTR7yZsrZL
morG7z+fBjWVL/4NVCDdBJm5braQU8+qvHUFkS2wqryehKb/EPn3UMpISifLybLw
mJEA8CSK7PYrrPRLB8pk8O5ZSTI/Rxb1Eayw1p5uQR/Qnzm0E9pm+RgNPu4diACP
lf8WTQl7JpmI5NIs0W6IbplUSjl0x4WNRuuMgTo+gGiSm/52ozBPEu/8n4Lwpdr9
LqLrK9zmTvMRlL80xdf2q5afzuCKJMhSnrqykIMZXvNjubF47vMhvaOGCHZ2AU6j
tqZvUUul9izPKYbqn3Oj/j0UaNw9U4H9Eqv6KTV9o+VPRnIfn8Xq3esAUW4swF3s
4TGK3iGqaC3dXgMVo47t02oES594Kx0pav/7kuJ6iZhC6FTN0hgkBZvUdX2JUWri
XhBqvWAIK08CulyU3vavWdyJ/Rmu0aieiL78yB/hZnNNKR6Nd7gXd/hzesvc6XP0
ijNoRiDR8KoYblkxlUaj8wxbBWICJ+xQ4R0E3FPFNyQePa7438yrbqPtIQBu1/3E
y4O7n1yvpDIfWNCZxWHPj6kiSWTfJdHrmqxZHSghoz5fv0a3bN+O5SEH6IbbYwOq
wcXcVSIS8UFiLv941aF8UXHUZkm6Xe/Xxt3PJH7InTAq10FiU7k39rKY5204hVzG
OdrTswVl6rOe/xIbtkylMsugSAMdtKBk4Pd1wXT77Bn5co55c3ZAqDIJxsuobeUM
iHRRXO8ynrjnOKB/wpCYLCUQe+X/6Cb6OCXXSJzfqQgrcbVe0TJwdOs4wwB5G9Wb
5qiZQ3YWMZyslAvF84OmVY09jYoyH1pYBGwbJZoRvbeWIrbmr5OxVpslK6KgIGmq
rtDy1q8MEkhv1VvzNNiYDG5JCvgiEgETgknPDs6fvEYEy60oaaUr7SO7A+34+ldL
S7pgDGlqhhOqwMQChcMEn7Vpwdor1R3P1r8XocO+LWDj4d0JQFhjjtDGl/stVY+I
SldHTltK4UCjOgaowAF2quNNb+veSnpPRR0dtJr41cgsqC9xMxtHvgW4Zenhb6ed
x/+3VEDmB/2fdTBxI92jdaqnoMGn24OpJuVAkBI5n128NeiY0rKTI+ThT1KElpP1
R6AtmgMNL7gpkFi8D0IppQXLXsnMgqRQ7Co3ddSoVoLjG9fzS8xzVWG9ho7G9UW+
HD8rRyVVj2pIiIBC5iJchu7lwuW1IV0BEXq/Jrkc/D81IC5MSAymqUt1Ag9XNb0/
dl18PnIMlN9x7eKnnITs8JaBCMlzW+ytDfphu6dFoSAI4h6+oTWS36mmJovlcepO
9VHm/IpO+lLF5XyO47lvqpLBL2Ouymvj174EdGe2axyEnicyrIk712jkkDaeU7Uf
wLxAZIZTPCuOnV578x1V1XxmKR94UAHrHS0j4R9IPzUaYZbMhFYRxUQYYfyu3DY3
RCldaNMLNlLXl1X421h+u3IPALZ+04dVXoUEi+SmX5c4k66wAa5VeaxamK5tKqJT
BGlcLhaUb5+THDXlIbLQ2uwHmPhAedIzHWr86sQMgRXk032VU1VQ7pyiI6xtn1ys
dNF/N2XVEeyb72R1bdXkY0DaktlzJzjErb+emTsOIyaj3VNFGyI1KhB8N06c0n7b
ex13//BGmebQoYfcXNd6xeDPKZL9Q4w+9UK9+JMWIiu3zAbvZuFYy6ZK4KEzu6Ll
di2/AjIquNr0vM8fStHH2bK90ku2aktoJM9XPRj8VF8m1nEpJ6iv4Jmqz55lOWNn
pXO2s70vSbPqpxiEetBNXiknUnBzz5Ryk3Gl6e8S9GCEhC2zpE/tJJjZJe7GZCOI
VBvP974Y76jDC2JAQvOxYzOjTIdYhVe6pTnIyVbPMpXtY6rtUC//3SSEaze4Ozg9
McccYkT6KtXVkoTimgQOeRGmEd7QoRY/rr4mxijRXCbNM52kSSFNt7aIw9Z1tTqI
X/dcKP7wyfmr6X+5GjTjMdv57TpZ093HoXHHm/RKamnh7TmFJZipeywBwBGhTJIV
jmcHG6dEhU4fHH7b/rn0q4mLOP9pFsE3Yy6WGxYOcv/fa+IiIPvXQs/Mhb48PF6j
vfqOAeI/AxScXByGTpMa3NX2GHYsDRG/KGsSpoUmF9a2Ne0lKdj89B+w2vXcU/gs
JMzesnd5Pny3RWQDW5cC4qIHDjzE7YYWv84GCDEutEYsHFdgCE1Q81TsD9oO3gMm
RbIhyH0njStXeFgWJp9xrSvjD2Dis/nj1VElugKDZU35GZ8FUahNxe0F6pJ3xjDK
iEbZ9EFgpjUWuo0LUKgoG5cTDToKcuM5VECctOUuY88cHJw+DH1f19YgMR5P6fve
c6ql8w37oTOqDeeO4XjgcnSHfqK++qi1NhtYGmc9iqFli8qgB2aBqAm7YxFuIGx5
7BX4r5wqTPyhtdF5S0ddYkX7SK0H3nIxXzYHkG7NQzrlacFHQxw5SGel0BBVyJQ5
COAZAi1aTzWFPYXuk5hCL7dhpjrx2OA/Pi73PAvVGqq9iGZIATMJxmNWzy0Id73p
lLTZor6mziDiw2laiblBoQIxwUD/VzYJx+ikSiWcxSWVGQbXOWQ7v401j/cB/bki
DSEZPTjjOD/dzmSQu3R3actzUc/+EmOVNOdZXN/+ALTjlo+A3xZN5MeUxCkmGFSV
+EdlpkhUcHGy3SETNcI5oTtCgJGHqacb269RM8+P1RIaC+M8zWpwyMMT6PoCJkgG
aIoc3nC+6XDHVB+zSCj8wHEM1p7trvMofngwe5CMIdnvewHk9GfXA8EThzNu9JhA
tV1m37RP1Txv7X0lUMNNabu7TF/XuSn0u27yHPDoKSMIKRZBOlWsTRTuCYLL3g5t
yjOK9nl6A/BlCjvVJb8C0F/1W5QtGXR2S4gKnPSVwegxRW9UnB9O9JJ4AnWgnieJ
yMd75Az/ucKYeyWUIEPg59dHDHuqAOeY+yAzojrEjgbggrt/7aOySdE7fUj/CjxW
UqW1z4XXutLY+HcJdLQOl1oCZ4nH4M1Kpi+E/73huUJYtJTr+jJT4r0n6qc2rlkN
CQNmnzHkwe3tJdl1shx1Uf47EqeRlx5qnRwfY08eOMD7n44n52iRPB6SIg4hPnMO
MeLpNXrJRS+S5DzIUpV2XwUpwcK2rPXfINIm+Q9t9kPmUBeeGyMOjQnOOCzw8bYf
Nz8W7Ep79efm7SROPGZXXo1qwgFqs6mqdQ6hfHw1hUuPLhcaQNx6VAUsiX2lqtaZ
BRii0TaThr320cI7XTvF9g5c3XJbP7NkQc8Zm3bXr7n+XsQYRhr6hjnS1RgZ3pdL
T/8MrtB8ayWgIuUrzylD93zmfEKXF2X65a2Zw2bQuEsXXwCdD07IDYQ91NheAoXM
t/C/b92uw1HBPrTwrIBs64K2kdIBAoqR5M5Alw4xYcsB864WzqoIqxAoYvmZ/Bne
xRfcAe/VFvo+14mTBbilpPSQWMyL3/v4aPvIDqPxfS2T++9xvQGyWFSfTqezXV9j
ogXGxIYq/BB6HmI6odBmwvukGA/+IPMcRJO6uc4Ll5WhWHwHOEX2/P2Cya+W/yt7
7jJPUPg8AuztdqrZOnld6LKNxZiVoT+EzzkUKUG0pW6Rab4qbFcrm30/TZQdcjkZ
PXy9C0hO9NBqjWZP/GAy9cgKzguM5iuj08bZEmgb0n9Ugvj7FpyLlnPdIEtCDKyc
oWrXgTj/G4XmqrZOCW6f/vqXDnyrGINJ8n6LvBYSnO8dfxGQp6oi9OKWtmpSXQsS
0GTltPhlfvdaZ8NWpzO9cLauDzZ5cUo3nedS1sjYp7eqpzbwyvqjdR70tVU38HDq
o/NY8nQve6Z+M9mV7sl5lcLeTsOH9kynx5gxd7CGtuhXPK8OkErPfefOLXPrl8zm
+Fmob/6mu8MYFrqRrwWYA5w02Q6p/nKmfJkB4PyW8WIF5zvd+GruGRTvckbNt2gI
EAHZvlHfG6rf+Q5Xi2ddZFlaq+93qWrmc4TYYQtAds3zzrcP6T3TFQGTDpdzP/SC
pN92Ss55bnY39AJVc9Gkfm2u4DzSxZekwTYdrddQ7BfwC7lmnMz5W4bCph8ggN+p
WZOYag8Z8u5B5UF03sFnoYjVMpELByRostL01rwoz7T44RpwO8bidddVckF+7de1
uRQQEEnwogMTz2eEjwfnPM3h75Pc/esX9dGp6q4uLK/ZbZ8vjHlZvYGToEBXd/+i
fygyRzlaY0XHLQ/XqP0F4mbfjAg9BLV/K5jhhgdoe/I52mPAOkl0MePyLCGjvprQ
fkxdzjqR7eDVVqBp3hPYJWkBnu8pEqOVkB9pTlT/LnLS1CQVC+OlFbfkhc4DK3YM
W8YkqTzIauIev4rrX+DWNUEVaF8jn4IbTg7GfOCozqQoCPs5RCOii+5ycFSWv5jm
D4H1BkSq9oGRZsjG5nPs7g2FnkQ8wL2sBtoGY33Mz0nI29xnNA7o2s3smKQ8KxmV
jx/dNMFLzDoJ8egiBvCDacy2hfPGBivEr9DXMHdT3UzqR5yQRXPajYq55WKh/pT3
I8syV1u0cxPxWhss1do7SCOqKl+jyTMab1Am+xiNuS3n9szrQkO/zLElEUBxszf7
twtQe0mNW2E21votw0Oz3T7XjXrYy3PNcLJBCyqYxj93iEZDpLF5IcXWCyzn1wmQ
8iC9IdkHFppQTzx9ktccHU+pUPhwN/NRiLZ3tAlLhBJTdX9gzQzZVzl5SFUg73AM
fMzRj3CKOzyVUttbz4wgC56f8+hA1gGlfIvc2RX7FYDUAw3r5SEmGKcYUmkM0YA8
Zund5UvRcHzH9/sHR4WZtzEDyb1Kx+df+YdDsZAhT8zYSy3ZQPzDkXqqwcR6FiXY
ZU8Q3TabHzdvw5iEswM9naSZJaf+zUGWXjUyfmmRY0OenZirPredwh1+XnUpv9Va
z9bi+JJ9PEJ83qT/YL15eKFeuDZMhKl+0oI4S6ikyNL32yqWLMjY/VBDQ28FCbgw
A2SmpeQyAb9scXTXdCGC6X8Lud5EHhGTHo+A2eGtJinLEo4qhUNGPS+cRjGJvlex
ltRyTyVKpbpFbUiAOg9KpXTRK1h+ccGQcTM1mHULmRyWCeJkSApaCjLRosiNg1bK
ju7KWjOm9qa63PZ+gtdJAeomgH/hkrLa/R/7GZMqvXJJ+BOn4592Zca4eAMxGd+Q
mWjB+oO+1Sbvoaq5LMCFgiUBJTDzQb2LrLvDFtEPGYq/N6QJfxoYjhW4cffBLHel
HozvRiFRzDxAKlNMR+2W+9jepqzxH1qW6hud5hgYcvl0701JteyEa4ge3e+0bf6g
8IEJeFtrje9f8sOJQnVQsPrsQKDEOZxjNSfn85SsYxI7mS6jJbGc4d21R3qIv0i9
+TrjkYPlsID1K2FMRC3iH5k+heGfS1P4u8yPIy1pPeXG20fwSUeqbyEwj6xXiMKt
cPiZDwnbQHeKAxXV95zkkJEf4pkjVx5tj7FuiK5NCJkIkxB5i0Wt8NIxHgDWXbXQ
pc9JaACKqWnsV8+daV3M+PpQmgOhKuk77RpxBdNlPGVEmIllPJH7WDwRfb0oXHUx
yZmvfd4mDQopaQCXk8gzPGXyzUYdmF6ufDb3S/DW8ymOPngOlXLa6BunI6GW1iCg
J9MZ2mgQ7ORsQi2G/05aJLKwGh5+RmiyQrYEgNQdVkz0S5c0i0sw1unNwQtu/LOn
0Nihm8cHktLrfPYJrjE688N9e1DeRfFjTuucFGpBmLK8t/mToifxI4L40V4bpCTB
gKdTNZsC3OAn/KOZoDd2fGHytqajCBcVZT1cBHrZZYny9DOPjaZSkr0/Xu3q4DbM
GRNCKiGySBpnAepby9kL/eELmTKvQ00PhOTRdInx082ECVscPD3K3tUQMhhniAjV
pw9lKIzHBF6+Dbduui4w6HUf0fql9awCxXTi8dfioZbsK/QGC9bU9ORUjFCY+d7/
GZ1DcGcEbLBqI8ATUZp4Ds9qR+mZ508boNfb06bkcqjLBf9LRotNGXvFOtRGfqcs
ZNf7zLqxspZnAAHqv9WoafqnSUL04qzkNGMJ7eEcpMbieZQ6UDggUzcnvpL5+pyc
SGQltwLHb4Sx3KXj8ALrFBbAk1VAmD+8WX9uKPhtuQp48HOKFO+UHcAuLCno1Ewf
Q1MmDLxTww76LLWg9sWXGkVBLJG084uS0Hx+zYXP3ik/Br5/6Ydr7QqF5KEDs9Aq
cze/1i2c3ahVTzhNCb8CuD6DCemPa5SkFPLkgg3chNMXng9mamx2LEvxd4UEzFlf
5qLue+5LZmHCpYYbR5BHO8f4M6jW185SSXf1hrQpPHdM9ch/CaUWFwdEM25SREPl
huyj7sBZSdYaiY3hLPfS5Soxjl+5NN8FpzZG8n1K4KAb3zixIbwe8Tx2XUEkjXV/
rUji3F6i7bBzbYL3LftzeasbhkpgQYKqdvjEDsW2e519JmNqPzPt9rJY1U78lwu8
RYQFXB8sAfo/pU7h6b+SHZz4xKrDCAIxclczTsNvEKxrxs41CO/9oP2UWsCBCNhj
r+EMXVeUh/8Lr6gYicW7Dvn5jxKXRcule8oKNw6nd4keopuLvJck6/Zpdw13xAsU
vxDxFkN+AcnUsvkzMxzjbqrpsNIOwIizbx7Lgj1b8TGOW63CvRIvSu21M/yGrt/e
FdYCe79qtJ29/IOntiW54VrHNj07qkN4zrW5vzbKlUQjcB/j1rl8icSY3DjUtHii
uPxZql4KehpSZ4XvIuZvuOTNiTbq/ZH4NqLptH1x/jNkkSNDqjAchuEer1lOVlFl
uc2psVigwb/FOf/fZ9vzxmcJ9XLabXsDN/aqZhVIZIVmTNTVTLnLuAzveM2MOgG7
IDI99JM3G78P4Gur9dNmDf54+VL86Nq0vP67pWCfWU87y3ADy656wt/KoGUoz2fU
U6pXrXBajNo+6xNho9jxTJJsdcLV45rJ2OU8Rw1sK3LtAHT36nVYgxp21abqElRG
Tr5gb9kfVtmsq1Kxw+8xqdzsNTOv4NyGLC+bOjZ7Kz/jAQwU6qHxjmK9F+gQURZr
HAbDA64uKs/x8ni7/Hf0agnz2eTIxsv9MA9zK1iqntANKM/fb5q38N38VcukwaQn
/umtkeuOrd6WSyXbNi02xFng/tGFcHH7qfsuQ2QWtjnaDhWc+ESttFzlpufThs3g
Yzz7ElS6VK0P40N9mXe9+RKD59PVg/BeZANZSkz4GhZrhqotct4c3vq40w3jqxLX
RdaywAF0gXwiuhf6EdV18GDxivf/YqPaAGqVWqdarRy87Wt2nib1BrWFz6zlRjme
F3Q10i6lm5V42fQ7yDbl8RgnurQTpBEP5R5a7PzSjlFspEhWnlT/WIv3My3UhUqs
o5RE0FIK2rwt4wWBUbkamCaMhRFz42SqXSxSMsiFAYyFw2IIlKvCuD+JT1yc91Ap
rKlKejViXRq//ivSaB1iShEf3u6OeZGGcItY62aQZIJidvSm8oavYhwbdKpyrRtK
kKO81aw4XcSA48wVH895gR737gcYANf072gZah4neJ7iZEeVUVTEt9Rd8zSxgDA+
u+6+O2P5yIrK6285sJ/TijQ83JnfxjEF0lYmP481xlYTDuozr+FzOAliU4BhPYPC
N0gdKgxq+skTV2FP+qz2/FH3OD532WcA5vV2zRYSxrTSQSR11r9qmH0qKUwWym5d
xK5G1I556XIS5PLDpHRAaDTS0wxukyVz9NhDLcWN/vgABYPlfSYxaOmx8iS0HGwv
Jfc8V3pVBpt35/ANzb6sQoHM4cLeAhLHKWoAxMugQuWMDvyBg8fy4/cOzsd7Wqtn
7s5w6o9bS6U/nOV9nTS9zOxNYyEBVk/2B0lYEqxsY2rpkDvSsdeOxVXUpvpB12kp
EnbLklaIEOljE6r+k1kUSNA2WFmfaE2vv3XU+QW1rp6us/Kn9VnGq4pjCiW/yAnU
8kxyDG87WtyhUMgiVjCdH6HVqyE70s2/QW5O0e4+9ndlaWR2FkdZNGjGNqYgbNt4
YUtIUhUgVnuiAvhERnPnFPI89VjFQiYw/8gzXEefo4Pi2HFJEBmm72hUKdXNGKxA
PfeTxyRfFUMxoqxyhgmdDc2e9pEPl9XhWVWqOHtbtIGWVkc2We71uZHIsUctcy6y
DFTc/hjwJ9CXtbnmKqjayhvNWNATTHzY5BbQTLLwzfu+Z3lOOC/p8Q4NGojIeQv3
RoTaiVHDOXWc9y0RDyAfnyM2JeqUWRZirI6TZLbhqkjaWvG6D2Ikr4QZ0uZFa83N
d1dtXCMLvOQMe5gThBfFz8jIQN7A9HCAywFso3eaLAicOgHuoTyAg6nyhHisM4he
erS4ktzPj3dHa9XvOzZDmmtoyoOfAaELW0yTI0YPbwEDD+meqmeQIPOaB11+bzR6
kc5YyhXL8C/m+mLLCuaC+b0g4UxdeY2TTjaqXyKMNgJdsEnprh2pjOJ2dmcWflUw
nAE7+Cs2WXEw3ZPQnctO1zzAx8UnxOfKgvUNOTwMK3UxZzyjIKWxJixN5bYfnMtk
Kt62H3879x0G5h8zhrR6WR0R93b3KbBo9q0KKflzhJtkaVf3e8OPK+pPu4BwfhBK
fj/dk/2L3apPxMTiTOcFaOfPELElX5b3FSqwTqCXDmSgDEayRvNd9maDHM3U3QaR
b6xXjUdp1iYViVz7fCukyHslDAYxTpWTUG7PQkU73QTemYKX0klWnfPyZqXo/PoU
dUhYB4TzQVRmQebG4bJVFZhSfA+VQ4tYwTibPBjHY/f9DJv3ugPSy/CFjS+IPFCd
SpG0+dwu13lbP2Ws3JEs6F5uyEIXukQIlCn0VjykS9MJ7kbDycWd47lBif/AQZ0t
8VDT+yO0DnFV2rqMmdepGs6aNYWg4UWuE/I/Xn1MVSTF6l5dwWC/sUkh7MvYqscS
lOA4PrtZw9jvsQtXqhPxr5SgZxd32JmibxwDWw+P2xZ0KuLYpa6pR82i5mhBbj+F
PLX5Ge8sPzYzQR3y0wIfDvmr7a/P6nYf/ySBccOj990igMEAjkT9dN98Zc+4xcuV
4PlQIChIe0+tTMAdtiPeXSf8yupEZipmwsdCbdhyBGFwIprW4wAbjh3pFhGhhfTI
d4gjbKsGXc3TRT9koffkQBY/qG5Kl4lLfEWV8pec+rDatydtePPnlKByuYLVzT+7
NesLtUm8u0XXBbzGyDvJ9vR/khvqhicVnWUhyxFYT3P5ptqTvaN2sz9iGYZI2sXW
MbmbNSB2kVg9tzmere99U+tdho9Dj1UyzHYw7wt/Z8k6jXpn8tTGLPpr14FybX0d
IGPsycMJLkbS5PX9nHRkR/iy6wgNEXFkhR1z9K5MtPSyQU1nnJjwXTN0odWd52zK
03mVCMu4H6aelgMp9N/pwr2Wlfw5bNG+0jEiC7jlJSUZy93isMYXzkUMSUci1ZYN
9bxyADA8LQFQ5axkVgNEm7DFp87KXz/vSRc0jka2NZ1vNDP/LDV9SudoMWApIWfy
tdgaaTM9jeNYzE6Tzxk/Nsxjp46pElUOmrJjMzfiQy7OWUXHpGqo/kseqA2PasT5
ke2olhXthKyCtQXmNJ9/0nebZiohGwKL0dT8jn6n+Ot0zop3RvskOEM7dJizftkl
lVRbGjuYToA+i+8rm3f2N/jU5YAbtHinzyb2j9CkFhDT1cNsOXdGzTtUGZfokhqv
S9TIWQD36tv4JQaBynoDTGAcoQ62ly3I39VgigFQ8ZNonypefOalyf67B6V4Co28
mi48VfGzq/QUddeZwKuYXPdnbaRct6+CsNnqPtZPitNARwz9yaBPDxnurbbXTlUP
M//oAptRxLT/yQQsB+dKGhgstYv1WEXuSKQGXiN/Lq3BClli+cunWtGL0sw4GaUO
BFbJX2tMtumFKgtTpH5vUFu4y+6GirCsIiikrIHaFOSuFMuRlYqXBgSx/RZqDQQg
FbWlkSRPoo7rlbEL7kGSjzxwk7+2SsOlT3TWTR/L8Kb7mdwQyySvu30/g7ZaRW4G
wGhl17Jm3CtZUgEQ2YZo2nQ45XL2xf35Kp6jGN3cHT5fFIZkMeKfN3R6eSOqCJhV
DP5L8X/dWaDX72GOfIoQoAW57QlGcQNrAK/HfIY+rY96VjHDIDxrhpMUJuTjr/nT
1nQmwPyG5USOq7N7EZBhRctBq7gN1chCR3lDJGRkPWVCHQbOFKaYGjUhrdCrLQxa
MbpE5DPWWtVoh9MS/8Yf8q6rRYVFcCcvQqMhnzsVUxVOatvB9peFpo8QKSpiNsIi
5w1rTchzL9jHgmVOUU6LVcrjH8dEhMX76WDMyhKPzakDOcRHXxDhz/xtaNGKNsHi
qcV8CFVEaHA2HvWVmjqNrJwiWjARvKyex/KaL6n/mZQyfJGZCVuj1YG7ECQPt5S3
PSkSFRPt+SbxzRamw/TUyj3IfagNpmkjeStCUxGpgB9FUoxMbyAYJGB8reHw91Jo
H0YuNzi3mTo9pVlbQlmyw7CCwhsa6+atFDPJay8+0DfMuwrWWr5OoY/NTjojZixQ
6YGbjSY4V6S034FsKAUuQGtUr9uINulS9C2n63dzkpvXgtcL5G5qX8GGiiEBdeaA
8TpURqPc4jpFCvfZ0AhU71viQ+9QdyzaKnzGeyFCV2FcIQDVgQXYVK9k+DZgJ9zR
8Vys5AGQc/RN9mHNYID3MeGc51K1Uw3CyINhxp2Hx4CHH0VLgufE/fw5X6PGTAkU
uqYpXNvG68W+AHWE3IsYk6qzzBKceQHiVrzmymWWYXqmzmnisJed/I+/eT6YoGLC
s05VVepAlRCcHr0jffwiL0V+MxrXEwyRFtyqfgyRbLT5BXJzBymJiKOnk3pXA0Tl
JBlZ3ydVtqVHaWmoA6FKUVMz5tkjmAN6+erVY5cdjr6zo+P2JxLOEnVdFkXGi/gw
cWRm1GNSMP2QYcAextVMMyN/eqvCf63zYxcxZMJq42SFY2GjPgZXyDbtq7N7tSMO
rSoSxw7JmEmyZcejUnJ4vzYP/48rVidv48v0vjKBkwXLpIxWbo93XChPLiaBm5Md
trBKUrf+ZYOi5ySBa2HDMt75OZxxr2NLD5OYOuU2qhQc/DSwoApgppgurDKHKWIb
2v84rHl6gAvVourQPU8FmK2bFVTBlObZAd3ESBu5tuf0j9iugsrzrfmwWQlMHBTl
WjPTQY28+J8KSrFH2R8nkfbUxQskJSaBLxVT62mMhS90ouAnuLvbp0ZzkfojfBcD
jxY+bQBcI/+ukoePAUJrtSkJY5WGslYoWb/oOSDMWIuTvB5qm2zjiCPTs1V+fd67
uaLHrJi09XeFOhnqrQtwgmAyleOB1D1O9GvzOcuMiXtpZ7/aM7mm5iP+3xXGtQjS
38arHVPo6jY+H5DfoCnz2wUlQ73pgwzQQpSKKzYThoJ2mJ9oyJuewIjes8733/jv
Eq3HYyLBgdYMvqRt/sdPSatHmhNynUClcruwvesicoPkS2CncCUauVsn/bthMhZX
0b9PtHUT7D19IaW4Qb4zHI9oylpVNsnixbANN/VkUxhcGrzLQdCMeT8zIq0BEyAw
/RQuKurXi8o1o2lN/bMbGN8LRssCcjO+eZ/GlJxol/4Flhbz65/BZMD5m+ZOyeoA
1i6mvyk7AZy/jXsqiy/GWy9Nu95n2VkM+ZpnTbVqNCSHTcNos3E162wvBmejZAp0
B2lHqZ8bVMPlGUi5n2LNVJ5QsQIizzV75VdSu3LVD2LXAnkq0g4XR+M1G8K7E3b+
AnNVm6+JJGPDwfgWEORnCAdJ9kzzsUkGVvzoFfZyf15ZiPP/OEENDT8wuh6GMYST
jYcRcLGBSyeW2vnTD+b3XTWwWTFM0u1eOv65KSLmv9CedOOxqhG90LmyWWqj8L4b
siTzNCZyumYyQw5Fvzr+TQ2kEObIZ4q4gYTdgH42NyR3PsgsfFVLnafxW8tz5Ubl
j4/76hBq9wGZzgC9MzZ73g1zBGoHElEykm8ZC6zxuxp6D+TiAVGOnqu4QJYAMwe9
cLgE5RSgF4uIHZge0JVHcLDVZyeMKbmh0UVJs5COmcCYCjBr5avt4pafLqDHv1D7
TkCzCBoCmwsQDMNm9rZ0L4FORDj8ZJexS+misKOx1hI0e1ximhaJodxBv3Oq9SwA
q62zV7GeZ0g56UB0dzaVw5r/t606BYXCJ5BO0d9pracfCcLl49s8k6FlOwKa9sV1
eD1jSr304qVBvXPvzWXne8ozWOvuGXCEnbJvptD7Qs+7Pl6UJNA6mfJBEjOeXHdT
YGBv5P79EJU4BbqrJVgPiAyVqQGDj16icU6dvoNu7fxbiffbKpWCwpphQRmI2ItI
mPIDR9gbonk9cTdPEi6pOgsUQ9nIlOjWkKyCYpBVM9iL9z+4JhAzR7JtO5U0ib7u
kZX76aIxhEcEUc5DPPCzpDiBwCO8ZLVNUIry3mHchwwEMToiXsAkND3VTP4BAgbG
A0EdAPnDd9ijgGoyc5wB4t/LH+NbstwAQqYNCcXkfS046CJW7pNUpb5OrYCYR0eI
nSLgDDNllhbf88AAnbZforAkCeI1ATE4Wb/nPBxjtntVRldGi8FbIdmjYiMyFsLT
CWLawP6uKaXti7ZuklPf3oxwF0/A9QbB5cJKA9cPZ6ocYq96PZ6PNioUi2vEmXsv
WiwxAGKhbVJAHjLSZL/GBq4IESn5O7/qNSNWoyaOPch+H6qGNXdZGMlLdAaaSVpC
tdOvGmjD72x5srk1YJwBe+3+VhUdfYHloRvD+PnKUCReVl2yKE5Dd0bXHhfHxTK8
vhRhSLi5zjBokkCYDQEm1V4vcGlDa9vyrqnANscMXQy0GQGRIu+lG/kRnEXTyZFB
e0xQGRrfnvxVtZPi8THNXQG7P4mIMUid3PELgZHxQ83lRhV9Jzw3D2ku9+ZIGVD2
sa0gQe1666SfKsGTLHqI637w8NoY1U6oPqsK1tnZEX+MO75omw9qlUKhnJ3oMRZz
X/Lo1gDNQYraRPpCurz/sljFRy95qn5WEWnxid5lkDoniuzKgnw5g8oy3Q9f9lFj
uKNgciOiEPi2rFtt//Unf2z9MOXL6+miW/TQecv0o8DlDvtF9QbuamD2F8iAJLHc
WqiCEWA5tKVFfaRT15v17dXpUKZVmuiG9cluilCaOZNS8wBz+JGZDXMIfMjow4FO
yQpzJrEPIS/moYC1VGExpUYMbVTvVMJVEqvruYu10T9G2l3rf4LPnqXbviTvG+wF
C2YV+a39uEC5QbDxVfoz7ycCtmpktuqOa18bPI8bC+qHZ+dwCfJFOIL6gVAUqUL0
cUQAIIRqE2p5FsdIQz/xdAaG0qt34gnJ4etryqRBzb11M39w/LuhednnUWyym5lF
Nb4mQ0GJzm30eZECVcG7A7ZmVWvAsAP5OnDw2g8I3RgTg7gTUN5yU1sesrXkGHnO
/Uqhi0LgOckgmea6XctvWJlVqzCXmu4V8xpu+mEdJDvn+bxi+DdR65uXalPXqgEf
O1hQiAc+Ki1+s/0U0UAf/jjgOV5K/tV4uLR6XrtwjzRZbHqw06yv+W3pjoOFiVfr
Ggc4DTtJqjN/xtdh8FjUnLpJVIsRG8R5JJlZ59iak/7vz32/JJzc6Xf4nEl/pQWt
Yf2hq4DeTJTxgx7MGnuEqeHNnrtXQ6EGDQmabMrIVl5IwXqe+Rf0xqTLP45Jsva0
FRXlOP/B1hLHJOR4EeI2CxaZgiK7JnmNdrBLkrVBybTgNqu4mUUQznY6YBAMmrpd
NWKY76zqOL3Prd1gYAZRaGoMloOprszQ3VCjmoBa8IKpULXE+o1/HSdZ2ihUJduI
Mx5SWNk1iDqiAjAlCzw0SEdQrpEf8WjvJznu8pnAzfM8uYirmTd1nRNpOH58b/Np
G8sGTyqqI7gpM8TiFJz6VR6G9z+w8RmUmqxRMOF9zJ1DXze7KGHReO6I437Qn2DB
U+k+jF9fSAx4dYoFpbKR/FIV5g42FudiLZEsDuT84nfx7YPUJ+zwsjzYONcTyLLE
RE4/uRxClhhapNdLlunJ92oawFsZ6d2IfxkgNHZbrQwYJqG3DrLtf2csCPRUU63o
exuCxDK3Gn61EiVgaf9XY8Qp4SLho34DDlSe+JBucJ3tayGXKQkYdWPRZeLaqAwh
vWMXQ1gkoRVF7J+IZIrhT4T7TMBbYgp8gz6MK4xuWLJdHI6r2b1AzLurRhXyVPco
BQW1Xw6OHN2NBKa4ICO7xvyRLNyI/7sYuSvXyjFCROqDsnEGm+Y7WDTj/gSx54Wd
RsK25iQ9+tlaueB5Xl9v3nNPu81OTZ+PEDtX2Pj9Juc1Q/HvVaF/hgS68nHa80co
HOgJ0+MZdz6fXAgPB6qttx7MIHPMM9dcPpZYaQ459B3nsSAfZ0A16W/nXcmYMxBP
z7V8OGmCxyzCwW5OcMoxNVnGWWUG8EIBNJ3Zhy6z20B9NkzCQpkVbh0G1MOw1Aor
RB9AwXPrWfvG1mW+a9/tQsXGP9BCM5/F4S43cA7uWuRW3dHYHIaGC1CmGUWEdt7Q
I1pgNnfNICV0JBhFnulMQT6V9AOd402cXOYNwY6j5oy9sm5lREPJ7VGp9PGmJVSk
cRmvF+J7QJiyhzD88EK8AltvxkQYLqXru0+jMLUiRnjamBYBF/ztFZ4vMpd9rE3f
Hory12UHtR337SBak7aw2BeXXGr9N3AqUvPj6ryM3pQd6QCspSqoKcnSp9gS7Dic
U6UFa+YSpS/XP/olUuea4HdG2f9ttAR/vzE+lwg7fst+DFkmMii/jir0NQgbjNH4
JL90fA+ssLxto7srzW+f44R2yiy1gz+bffzv0pukypj5AVlucJJdqQib5utPJQCY
jO2ENJh7JErjPjxyI8yHd5Cpy9/D6idZtMVkK5CUu7xt0TEyvbyDtdV88BOH9j7q
EpXlaK3vSXnPGcTjtMJS4Rdo9Pxq/7cK4xrkj3uoA0pp0KmIVf+Vjl31A8aapwnq
s/iHS3HQS4IdXmk45ErWj0UWbG/WuMIFV9angebv4OzIuS7oCduTkAlsmNgWLp3i
FOHn4f0UB49OgBYiHkKlkRmptcvlhszJmQlEgnsCAljw/KAoGWXfahBmFfz4XXa8
VvCuZWW2538KVRZoHbhBMn0KxlN2MIugpZdvwdf8ImH+LgDEhaJQxxXZ9YjxiGuZ
g+vE2XMA5kpw5TfYHFm6GhHFziC+w6+8wEfDYzwQ3EVY2RWPMjlEP9UGNakeYLDj
TbOWpbFhnUUkTIVvVImofJ5dQyUCBzJeY4WFPpSwLY9xvk8H13UYZHNl3kBUzq46
xlsbq/V8emVr8BzoI3qZ6nlBRI9qnW31E2drDSwTS+1PGolSZkF/PJRaFfCEguZJ
qpzMlCGbE+j1mXaDtix14lfJQK74mLd2sQROmDzdSv+cACXuOj/bzLq575ZULGc7
8BF5jadmrrtg8NoVKsYLDcCJRRVNb8eHdjQK28MkNzRDwmFXtj5fuuqwnRAXrZxf
BdW5Jf1uDYW9ljJkQ0tQv1KU0wDOJ3ZFA3DXiF1JmMO9QQ0MNB4Y8fkp6ua4PDWA
ORnlnfGEJ6UUyODG7FI9YzLplZcaJnfyHb0qkqNIRu9hn8joQhMwBXpjlZ0DAcjb
m5TB0xSkd9M2nke9j3r20hlD5T5a3K+bdsuX3pdAJYBPlRikRZpCrbYzGH6Cj7p/
c0bUl1SO8x44bcm0fN/GrAYCqO1wwJJ/GVLKimUnE6Mjj4Ps2pgf5bbtJ9UU7MtU
J/t10q/S8mgCgY5P/Ka/8rEpSXEhWQEKHsYr2RfU5u4QcpYnm41afQ9SzMaICgtq
R4rUQu8acIMb4H7tcT6YFk6aLwB6sPIB3IHp8ED1vWoLCgI3Mi2DdOi91cQwFfh5
MldZhB8htHkTOf2mTmSeB/8rNGOnz260joBqQcAZ07heQVHzl0PFW/dQOAmDukm3
E3nje/KrA5+4Fpz0C9R1vBfWhFWPOmzeRRHxB/E9QhcQTz1Pijb9Z22OjfNrEABW
5dacXsTORiO4DGaczgCYHlCHpmySCeznj1RTLXhACdVynVuSwz/gtB7fvNfcdqjB
Kj4Tv9Cz+L8uilY449BHBxdoP2WkRAJkMDvkRhA+/gsadIKnhiVtD5/GVaVrXUOR
n0PWU8MZHYWtuv0PQpELLvOqgEWRDMK/tbcgrYD8rgauGtF9FwhO19ARJ6fjGuiJ
cifci+0sPp3sErtenCuuQYL7LEuNy9FHvoIZXwDcbX1b6e1NjazQ04Afo9Tpksm0
d/4185kPho0F1QcqYiYUnZm9cSD6/kxT8dAuEfX4xSxwixLzSNkXhdKaP26qieop
ZbZQlViqb/9cvAEhHb73jSiyda1vCRdiQPv82k3H5z9aHWgCc4KCeS6FbpOduin/
SFMID8flS0zb6W3ktAjs4ltoUSNvxdxl4AYG0FTfBKt/MtQshPYA4Lt33sra1P+Q
Tpx+SxkkU1z3/CscpMPpTBe7mudwNdoX7rVf3ZWmbAIGQC3I3VrEoyVZsDn5zpGO
uL9uaejQrsDHy0JFIBPreopequ703N+kQiaCfB60EdAoXrmMOnpzkzao20S3uhKo
AyMK3t7Y0v8HyDuzzXKE4XgIfxmattvoRNtkrpJpSaxmWlpVbjUk/wUUQjDJDGnm
KqT0uJ91H+sNiwWcxHDVjdzfsS+PUqmHkCn1rtkDGeuUi8uhKltVj6vN8ixmSnnK
uVUAu58zpraHk+LoqPRQE+S98BBR0C+YyMmu3p12WeDUu+HdP1Kh+/PVKmZPrT79
5kXYb3x0BmV68FDFgj/EsMXlhDJ1xlsCc9CXTZFwb358/7aLWY6+NBFne2ABTt4K
Bsb1MWYoC/ipIKRTSUAHiF/6rPgD7isLPsAn2prRQ1+BoOATz0gfGB3Mzx48XNUU
53mJGzpEPdOTQgLUzAjlenl8aVi4cyZjpHgnrtDXR+1AlpxrZS+wGkAmvvEdNKqA
LtUdsE6mCogT+3VAh8gbApelBbY0btW7PqSoZZJGBNfottxYGvlIeQzL8ClZpPON
fYaZ7Fi+KtOZvhtY8z8IlRjmz55CnozyJwg1oJAEvZ6g8pA46hl9+q5yTeVupcDv
gZNB704imwZQythxpWfoxhr2ruHoi2a4WYfoTIorlIlTlw8kqRWLi72mF41fxi0J
u/s04VDc1mHGCQ5Zg2APs36D/YYAUmI/RYNei5KQKwoZHJyOSuPQfGY3gXlwSIEo
+wMzpQ07Qpd+J6AE1oXzJiJw6JWPb7tuyD35vb9k0EiAJys5pBU+gJBSKq160vaV
uMHpIp7cbqWH6zPxoTKHtkUzrSLxOKzfdpqBWTv68EjvgcFcfgPKdajYx7DLMlg7
nfpmbatNN7ibDZWBRuD8gH90WwQ6CbpL95o/ihsV2rCP3sA0ZH1FFgqiXA/ZHHoS
YjY6uB95XTs5Dab0Aw5vc6OV7jp+Z8hA3wRJU8OVw+Q1bW+8e3xrpUM/CTGOC51E
exin7bZX30OgEKZqNrq4WTLZvRSvfoahxXGgUpY8XeFp9iTQ/X2MLR3XM9fe4UZG
ZT2m6ILmyjIXqU081OrGQSinyIIUJXMSi5n8ZQSc5tw6oG73p+fzYRPAgGEJrZ5v
ecYhMpLu68nNkBOIu4w6ncr6WIJDp8Jnd0IfCv6g1XwNCEv9g5q9PjWzV/QPB6XE
vq4WOzo5pIQzSNI45vA4kBEHxjTwrKe1nXS7uh1Ufi++anGmdTCU6TO0PdbnmQMW
wyogxjOCCoyIfB943FogjOS+WDY0OdbqxIlCIGX4wntYi9gBMF15HLuA79Kks8uF
E/cP+8LGJxiD4ooeJh4ZXHEC969gEISrIm/L/vZXERptIddL0kpoIi7H977y8svs
Llwu0OYiZPAfqyunTxw+qWYswEph7IMYzOUOsrjH33GgLn8G4aVJOVGcL8k1BMmU
+/bAvoTFIlxCMy70qH6yhwyoyvgSuaox/JhrwcbVgPIWh7HbPXS8oTQQwvQemjzJ
VMLNVDdEMs7OiJkAPXSETSG4k9klI75sa5qzi0jHl7NSHYqfJNiHsdzzQieQP5g0
7Q2wD7YtOc/ZqIncOhtxoEHfgArXT0L+DkUREC2bzG0CSEfQ8Cn1RWmrdp3V4jRz
yEi+utIMVlBcK0qxr+S3IKSsK1ek1GzTDNAb9Y8cpMJvj++YoElDRFNt+EAzj35x
00DUqD489uihcZGwL83PYS7gD+o0p1IM3WR1q2GCwnsqHEiq4AXKIQbUWZOG688g
uhrD36GE1yLNCcv2rLaizSgBbJoXFikkMiOC2TVbAorO/01in531sJV/ijFVl0Pb
zRJ5pUOx68k9gN7gOc2biqbyWMDt/gyy9pwqQV4mae76WE598bADZVwfoKq8LsIM
9LMkyB9p+2G0lfkzyhfz7xkdbRz0lffP0N0jBL21ZhSbCkpjzxOjBVhj9VvFTuFd
cN8ufPDv1nPEqdbQ4kc2IcIbvOdja/4lduTrjEU09sU7dhbTKjIdVzl6kS1VzWIe
l5rwYAb3yaUr5G3nAfl+0vz+ZlktrcRLUq8U4CcR6tROVpYzg8XVkIT0UmbqPcuo
XLMmRt/3bHY3GA9DzMhrwq44LIl9vVqukoAt5AifKHZ8HfDN0PyWLZpfqL1VGlJb
aRxdZA2h3dqYC7ex9S0Z9UkZXSshIZ3fo1eMpOmDATjuljyExNyAb9IPmZXYTimE
tp8i7tMQppE1LpGZrY5BneVYXq69uz48mHPgoxImI7ixasyJRzjatr6ppbCi/YLe
SVH/yLkYmqyTSO8+QqINrxlt7mTXHT0YJekOUHzK97hF0zQMPxrEb9Q0zR6v4v1Y
ruy9nOxexLzeF4SLSaZtbOSnahC6hrnl/vEepUuSE2SVUhRIxqyyGNu3TSCZzuLJ
SHuQ94SUB7lP53nwuQIFNZBIT+8cA/rWfpu0t2S7Ag8vQQsZxr4UnCQ8rFUOW09i
legVCgCHqh0hJBqR9x8Kzs/To/HQQ05S4i5Q+eLORidtg9EsbofIjAGY7QvJsZ7y
7wwHARei49mFrDRebim1Jw5BRIXKRyvlXk+fsm46ZHcgfOkLT73/CCBOrRaGqhLS
jG6wyEkf2bzNu1ce1xo5f6YgdLfON9Gejs0s/q/NGxfcm4Jq3CLR2lg7pLZ+fYWw
L1v+1gDcES0nXrVoMj8bEjEcpNflghJUA4CGvIRqKBqIS4pvR8dYwq1hgWEau/x1
/siuxGCBcPZvHtBQMDuZ+ZcMhDhZ/gr/Tjh3N3kaLhDpj08s6wG+IOnUWM7BvsLz
cqwnLtAY2YKsUrWgpTbkj/kyFf52nDGoD+J3KHdHaOgVoh9I/gV4YU2GrVqPg2Sk
TYNtY8Ovz8BfS8LlSAtfiVFIm3px96YaxDV7ue3zPBVutm3IVWVVL40tK2urQQKd
KNOiUJItVLy+aQhSaSWZQSiprx2ucE3On3c4ctV3pfJf8YCErLcC1vRG1QezvdlA
vRHza6vVlvbSP/mP82UofJ3qVooP3JXBKv8xUUwlUy0DlOgO1f6SUonf1nBQJnHY
rRPB9G43m1Os0uVrAAP7E3e0Wwkf3xFMv/xEh3L1zuSk1SChoOibEeJwU797sKlp
z9Wnit6sCRyHs1lmnQN0nEsoLjYWMA9KIZ+IutwrTAP8xXpXnhfDLe73OR64LCCu
vn/VkFUkrdUD9F9XqV+KwOZ6FWkZAPqwkMxS4R8KE3bJAZNGztkA4GoPFkHzGzQp
Qtbeavdg59thYM5pN2J+7ewtlo7VtfyZ++Qs+mYr6p4LgB+KPTpUJG1oIrv7n34w
xi9GxNRCbrIL9FH/3S8eNJAV+yzqhetS/ghDdtJzwkQPcxCYcq8r1OrtAoXTBYFv
+iSgVXr2IYP/Cd8LmLB+2Pcov2fwrVBNAX/ODzUghS2fQ9crwFKM9J7fYX6Bu1yl
mN2ast2TDMNLGA1Kwrt6rcW2d+8ZbrUt3rS+ftrQnNxWD30JSg+7TAunAzUQMTRj
PZSiKAEDjM70Ow2BXyI2luWmPHts+LcLgM77X9nrEkOd/CdgxzK4ahsvbcXvy7C3
dloA1QaIJgrN4rE7jJkTM3uTECjy1OTP9LIlFVnkFSiOHl0c9GkXF4utc4r/CFtS
i40J0FFLCdMbXSKL/HFrl6zhJYctqPmbIYS5IWH1wAGX/Qsn5H2Q68tW7LZiUNbL
OUvaOltTaYto44nKcBukjMWpax8qfjYtgDbNrzR+0Nv1BubN7fJ4MQ7er8mgePb6
aEdzmwFitxvfSTaF+Qh3HWJxaclkrMHuoAMgh9zcB+eEGBoASMM9vtFOWS9dTpLV
5veCKhIvyb8HOlEHkMSegU9nW+1avFmdDCrCv3G2JDi6dId01nwjfi3gMEpdKR8E
PXEMvsHkR9OpI1YS3UfgDJEY+PWq806ED9XPbBr0MrwJf451GGFyl4HwN8stG15L
ms0HhLgzkVJU5KQrwhTs1KVdeOjQEDFSBsFZg5hTEwPc5h6LP6AuluFkW2kvJdWQ
k3EmHuxQrcyVjGW4ytCnGiN0kKdSHNuWsELRMbqaR0KM3PJv388uPP2YVTlfRMuc
zkfYfq2mhO+ospLh5z2u5Zo9ZJMKD4C+cfyWfBO9Z4+2w6GuAdsO3pw/EcnwvkDT
VVMj9K+ESZ8sXqYOiKuMymmStKmNvVW+LP0mxsGUHJsPkRAJHQ5ERGF7+2ck/zng
SWH5r6vvvmRvwAWcQ2vQQhKWWDJyIcvoOrdRZuAah3rD3Tx/RfVUkK/2I+cY9HEx
Vd7f/4yxbi5BcxcWfbvP5CW2XsVbKxRYA4K4M1sXdET0VQ6DSSuIxqG6c5xHWAhk
HNQKZatgImHFgg7umZvdQnRtYhdH72dlmFXsa/4DrN7+U1snxS72u5pbgP+6HsgU
5n8Zukm4RKnusQAuae2gwffrxMXo0HvEz6WiYMvrigb74b10YtcVuoFTVExk1pux
fqydWph/yEe2weTxMBy5LPrxHFGeIy2HEHiB1J0CDWue8XyBMiTTPPltvyOeJuwN
od1m/w5Dg7C9L41bluOaceV/OZOhcsbRzK/ayoDon2FxcZOP1xYC2cE6bVpC24Br
JT3Y9w3Y0n19lTAPlmWTsH8pAR0A1IIfpfsPA5E2dsfQfCcCw3En44cV6KcxaS69
eLnLzDfP8rmunIR6dYYN4IQdphXTin3mFQcQKi2xVz7DDRH42wAcUKPj/H5cQfY4
ALlPTpI5SbtKyPJFn4UAYEKyhKocWf+lufVJLMjwrZMMvh0AMZ65oWj+j8qv3iRd
U5bXrIaS3DWYpuHlMs8Mpznhugxgc+l1KqdjR2FDUmClmkacmtyhVfN4Y1NfkUCr
jWT6aHwsQySKgH5VwCGA+RKoo8BRcC2Qu1oa0MQsnbRk3dr5USwGT+pbuPUPlEAD
qDL6Ro9f201TIYT4tj/kZW0udDU3eGh9SEAUyt8R9oE5aa7lqYXUQ6OCoJ34fZpw
FHtMfpdrclG/qcWZ9xpBe+dczjO8tSzk+0bZ9fs/JCxAegJor4fex8ViYcVSwGej
o+t86sgII51uzBM6YrXmfwPNhQNxwNN3L5fBn06mdjQuVB8tNIn0UWBZ8cXUtpzN
tE/HkQPqVLYMI0IaSrSsn1NxtInWRFeRS5Pf+HozrzZHGhGwsgIVg77sqEYgzWZU
O6XVCww4DZP8oQtsf+sWOhRQG9w8l9R0sB0HNKTrb4tYQH2arO6ErHszLnn6+03C
uLXc6O+/Ws2GcXG7zGQB5uvflAFEzW7tDpTyCOGI2/pEv5wit0mOt/By4Wg/BsVa
YGsLNedC74CefxdB48UUOgjSmNpdA6cilK9U4EP4ocA+3gqPkRtChh7Oms3Gt7ix
kymQdW4UVfV7fRhbjX0HwwpnxrLqoZRha9Tc+gbyc/CrSjEV0glG30zNrY9LEvlb
OjoPjHyXaBnR1hDj0xJrguLiTWYOaJIgeorV6VXJO1B+/rKZfL79yQ8/nzSMPbO7
n4sImc2JY7kQy4VJAhsTv49fDRMXmFmRnG2niU5yY52pTS3M9jGooL1H3ywwyrxW
LNxH90wPRPofWPJNbdo5BTTwGdHUa16bD4X/iL82xAbPwbUQW7HdDG8ZPe7Qxhae
AoqbPszBG0iyyJ4AzeELv8KjQkV1g08LXOAu8dHbJypaSFfLUP2g24csXCC5BhSN
TktFjG/sR2zb+ek8aVq1RQrqTEoE69P+HPPo3SXlQTR87YPhEEdXDWmIkY5yArgi
V7aolqmjU4cf3uM60xyYSWts4UuUgSvoInDwSavSrUoxiMgviuhDeohckpqm1ghj
mrNvBx9ou3plzer0MAL+Mjk7kDB5djlLWH8B2jxLLK523i98QIAd4wtsBB/Ah0Z4
nVIRASOJ1JguzLd3/6X8SlJU7MSeocf56ne3dG3ylnrQH6NyStejkvzQHlJZZdJa
LGpfbrNOiVJGTigjmwg/wBG0zrYI/qgsfxaPTijQQ9EUW5+o1l4AQE3xOqoC4kOT
RLSLoQzP6UzNSHlKJkQxeOzu9f5MlcGi0/ICxQkbhCGrfpZ/bphEfilB2eBya6Sz
yMW9VPYzP6ZlHggNkALbFJ3rLZjDb/cgeIgJ3UckHQi8E+s5iNXfymCh+V8KvG5J
wqpmnKIR0ZC4Tiwd/ZbKjVoJJNZdsrdUgCZlTrBAlRuwT0ywF5RaCj6ZANbZ+tbJ
fIds62QcVsz/nx7i0qR4XhiVj5WZvLgtPwB4MMRtVILYPFwZygL6ELnbpbuwiBkg
qBwI/ioWJ5oo0YsAKeVHy4J3RnN1GLsLoPwVPhPE7t3T+sqDgSQSyqEZBouE+ZdO
aafzw8acETyhzoIoZ7AiQh4jwkjJzh0YH/VzEkH5csTWQ/dnQRG8y3lZEo4T/UV4
3D5S/+Whud/d3jcGs7+1zj6OlcO3IHIzEPU3LO3uONEgm9PecNHsDS5r8oMFsnYG
sDeAV7d5jN22kZr5AZYbw3Pps5Vu312bnEFmy7c8EYUNP0S5LZZyW/Qaa2O5iiAI
mFmVsVa9Vm8WspQACsiuiEHodTJYjoiGTBJQnfE3LWDwKjmb7VBFqGlyFsEAiJsi
HDb62ilGWcS6/CzzLz/nVVRwe5lEjYNOQ+8enCPQO17DQLZjoShieY6jbMhOnMLd
2aKhoSDSS5TGGE9lNNgCTgycZfnRu10SVIs0AaB0RBXNloUSA6i1ERWpkSljRpY6
z5kwlhDdHkQyIWS7GAIW6M277RwUrUrzw+sCLXAlKgpBpH0PaEt/2YSYEvk0f/mQ
aSqieAiSJSxNSMXH8IO9crnLYYts3x2gt8otTAUM2d768m5QFr96IG7pbYprquvo
9tpbrYYXEPn1G3iUM0TZ8U1yOGuFFimqqbb6yIaIcIPz5d8PFMmx47TPEmScZwck
sU9Zumdmw8cO7L/eebjPoCoPvaliBP/1XdECZzgRtkmBHbbG/6Z9kajR58l1cdh8
4T0LeXrKFjgQwRJjPTK1tNQpYnDmU/ED8943gZbU6aFjR+SZUsNRv1sZ32fJl1tL
ljSV7DsQ4ujaqdkr4Y6EeQCBqcpcz5GnT+6wpgQ/ocVx3bCUAk6wyICemh4Mt+98
YNVbjJGM6pqHWz4uZmmUGBM8YSTwGJNkO/BSalqRNWLtkNQIDc6h3UdcJQ7jsloB
JBs4NcMxZEKyeRsjnfO8VGoykuJvS0TvSZ1fuCz9laXaWXqPFycFEJPKCdH7p6xY
bJmOCh/fYGxic/83ii5ztD+MZkG0L0MeADgNo3UgBQPu+tYx76cD5oBIMSF8eOik
WiwbJDu9OAmhKRLGatn0vS1gc7D+35nWTDR/hg47aMMS5dtHRmbFFzMSfSrYztch
VjhTis8tuzopQkmF3ki27QjX2mlZRyJOSFgW6aySeK763peKUIlMXrY73O4xHEun
6xXtfNtF84mUtMtIezxMFLXBvX/aYnMl40qw9o69lcMI24x1K1CYEy/7C0LgSE2Q
/6DoubMwhOkb7dOb9Rop3SA9OM1dgHNkViev905amjxhQmVadZYcBbBKr8wcNpdv
JX9q+1prKQfMUdQio8hNwRAh0dRI6lsgm+Rr15vaF5ke5xV57j0y4Fe3SNW4Fg01
h1C17gMqyqxne1eOHsQnpws+bBHLWbUdvzWOKqauo+n+oglOaDXCEF7Y76K4Pe5c
Kdm1gGxlzK7ySGMrVGU3e1tgqIHtlFi4djRuaDfY70vFmxpUTzmT7ftl8UsxZua0
8V+p3S5wCZIrx8OMe3ly282oJAgy10GEpnqoF3phXlv/TufL7ZtwlnZRGpj23USZ
TSMZuhwFDqFLMaho+v99YkB92njNKFgXPXOtLAPoQNznj2Q/MJUzgCuRJbPSGQHq
gm1KoNyIZ/HQ9B1ZeXeQYtG+q9J7wQ0nVrRozlNuvjlMK/w8I4/K8qiCulLn/kWM
/cA6QbTOvvgUmEJbTmLnt/UYy7t54UQd3uAgLI/qVszp9FQugcWczvZ7ZCUzkL8A
QMZOwnUCQ5uTn9vmb5fBgIZAM26Zne18o4btTfmV2xexy/2lZoJx2J1HndBpkZom
ZwX3uFjbI1fBHZ0KwOVEIfwyzdgrFf1UGhUmusZuqBPx8a/YDxYsCJYCPAQ7sUsq
kF4zXzglVCtByxtzBnCeF/ZwcBum4vDoFEn1Lf+f1oDc4XGM3sPWHcNRvNNfnUNo
Kr7uep4rcIP0M5lOorrEH0x2whaN0OXoIxcLQJuUOKPSqK8kp58w2lTuN95nAvDY
VKzHe0BzMU5m3DMZ3Vo4aSqZrW1UEfPRlEWvpdEFXEnOdc49nYM6yE/lsCikaS8n
P21MQBa4vKCyRuIaX+i+f5dMtcaDIGcYbzVoUbKY9V+RnasUMncDw7XWRlRAjgY4
7sQUvquLwAImSx22bIArgQjDemmbdAbkREI7Kkk2rr61uz7VqT36XgiC72VsbfKd
s2eGdUk3gEgjETeZrZU1x7D3adhpeaWa3eXOrIeadvZKRpb6GBVwN13l27sOLVmP
/5FVaa+tfE6gyj/pDdE+CcIljhuQ/1oKXvmxzo1AFT5z0VA2a5QLUvbDH5/YjHdJ
X1QodWZRT65gAiCmLLXrAklWLCT1S9V9Kzcy1nF1hZKT/CMwk9eLmN6MNNQ8voqB
+XiOwruV7ao31Uds9w2l15Dg3bnhYLEHmUYCA4EHjuh4uzs9jzJuIUiutxbEBRnh
h1j29gdUcod/Olj2paXR7CL4SkRYpHo4v9GdSAb8TNax8I/uMAtDaYhLp8z5Vmf5
BGT+25/EKO0Xv15uSTJ6lzl7XObDCenRivF7YnZLla+GZoGCZn5xevAj6ZEnvqeT
IXB/Tm8+6QyJstkst7YRWkUvNx1ZsPAIr1YjW8bVJzBAtiog9lOpyzif5Y5Xd+Bd
tY3MTbcnClQMQQg94owMbPg9gMoQXRP4hprjAft0qwcHtaXQDt7X+2J5fg4hu0Wp
k+MwN29q5yZAeTv8pprRFRZ7UUhJUsupVpUdJhBj1yydk4/xDPiJb8gJHjhRF4Wn
Q/SRVTeLSUQLs//cPNPnn/B3DLAF3Qzom32lrb4WfM5z6zs1ZrTZfkxiaHkadvsz
y2TU6JhOWzytBjXJPF8kzOWe4qMp3nK0KuhkHewGjH5NvHDY7nRSRzHbhfo4s14L
+0n6zX5bafH8Fcfsg2FfyKBiHtIivAEq/0C+78CrZUIekwXRMLxPv1GUW8gG65rX
Ful5E66AsmY3B/IxFDHjFWLXfz6vR6gHoL2mJDmSM4M6AMzSZi16b5C6hHYVASNT
YNebWgV5egRmdkngs/Qaf1NK4U9XT+Y4WXkO9SzTJKnwBmBAPmSnsxYqvRSOKYra
21eXhLB3nxzLP/kTkdMmE9jqrMZ2Oo8w5J04wycdpBZ36MIONftygiipY/0/0xEP
dlTB5dfX6MF+FwMa50AR5JtrOM0yMqPPclObLw5wg9lBaofTiLg1xdmJ7dObH4qF
HaUr3/ZDTz59BwQPC9n6Vm5M0SLAIF3Gutu24xKsguEmYloFs1s3nyN+e/KKXqL8
oIQz4rTah3OI7zAfOLx72r2nh/9KH5ajUy3lbbYtACSn0iTl/q6hJ9UyaM0rwpN6
Z/eCtAhQaliqTszPIQ3tLkSfz1WGLkZSFEPeSclMQQdfFag2UAqAZKsf6wCfTSW/
SVBDX5uKNsgokKjMBaqd/3RKvhBg6D1crfsP1j7ObWVsZ6yts3UDlwo9+2nP2xnw
CZjMerSLidSQ8dhFhBkchsv79Nc+bJdY+7z6lm58Mspx1QW6eNKbRmXnSQqwXr8p
hx+cifnToJzQj3gVo4UEA/AfpAEn/oeqocF7pE5ut2sr/hns650A4rOsU8CMpugZ
N/nz19hm0B3tF+oN2tjBd5VcI52alPn461oeHDdGZ4jieoTHObCw+mBwe+3/yqYF
v3vd1c8GHG12LqfEV4IT3WuGzQpWhBs7w/TJnJP9EhXmLiZ95eLLBX1xLsHYCY40
BW3CaS3jCi2mQoaSBrvAIpSy5wC0G88fTsQhRJUfmwTIL2O4+Daail1lHLoNEeHH
uvYcceorpIGzFlRqFzP4p6+ZMmiQMH+XinP+lWgZ88YsYsBt5+c3EdN2tQ7+4MLH
X/jsFp7uPo/yhPQlA/MtlLLicGuNDtfMeQr7/G7LBqesjJfgGjYjEju72m4iJWTn
bLHUn6FIusX5AIMMAhzmIf6bFYB9QwgHu87lL8rSkXlysJbxQWnULUefqWXgytHR
k13AoVaXv3o92GXnrTQvMRnimSY3xBH5sU027v41HU665QK3aX0CdwYt1jmBniv+
dYKH7sliHcMJ3El9F1MKZfBSvdDFOXbZTXLFzir3JW9ntjuinCmEQpUdncJ/4TQJ
tkpgsOmcRmQhI3/jd4quUQCu+u/5CJw5GW65jd9/xSYyRb9ecF8xf6RBS8pbh+fF
DeM7QArrBKPlfgwki9QmjeO4qairWKVd0jB+HO2+7s/MkcHSnicAKaGK80yVHCad
1hTlE7NYtXwNDEavZ5Ad5+szklrFXgE/ET10bOO8l3aSNoGd02eTvS0GX4l8k36K
oRt+4s3oCaBtaJnvUBz/4bjvqRlRg264q+FUz+4UIfsZYBbzYvpPau6yYksIA01L
d25OW8KiNRIEwfbibkJERQ2WBGJjVxMp1Ylf3sYOxw9Drz70HZRG0Xdt9Mhn0CEs
t2TX/gdwJEpUsvpU5YW+R7KEOvdT39qvlxnDqgEM772dvQEhNX4f8iNiXGLE4lCc
1hb22WLEPymmld1rt4J6wMDfi9buPjzjLU3VRK0EOgc3j6XW7nEaPBjgmERwQ4dM
RlueOX+nzIkWybF0oogyrVUpZPncvjW5iNTHqfUO//ryEmvxM45dsCBuAesPIZ4/
IOR7RRbnrwDIXHVJJw7flhIW6z4j0IyeODL2+mCnynRVwB4VEh0x5utsG/cIUbsl
uVv1uAZdpbB0XXaJmTb4m55ODahymrXM0GwKSgYy9cKuRD+AViNqeMh3YAvgF5rQ
EYsVxMNb0KNfiOmARMebVmA5o7JyX4FtWdMQ1BfARZ7pmLIPlv4IBNdmU3vhUfvS
KlOoFECk7Q08xyo6t/1lbs5VHRmwxHDsF/Mlqj5ntRxNIH+Sz2/xSmhu8+nzT5eG
DsJf8lUcLRTB35+aEFTZwnZgY+rVr+RTfj8ogyPI2TSNWzb/HAPPGa/TUcXZRNIs
YEGgaboidiHV4vy8DeQBotduH1S+26nexkYF3AvHT/AkD/t0pSFkVX6EZOE74rmF
VG5368NAgEm/tuXXHbAbRZe5yf7RogR08MZanUYRlSMeEqRFVzNpkbSZXvDy7+MC
VrjvssJ03IAesq9kK9iy8XlQXntsYvYPbJD/a4lQHdCCrFSWhJoSGdiwsCU6YKbZ
1wpexEP+Mb6lz+LPUVdSXsTlLTYcz9WPLuSl4/CuoWt/ltUweyilYA2DQfeajqzo
ZwalVnE1Vk/rGAC3L5nzijWO4WR+x/5G7h40felRfWAzSXXDeCqF0Vks/K7WyWLC
hLcT0gFHnXvujVPqrgYM4WQj7Yxtev5pngDdBKhHlsHrmZjFmiIyyknofAD8/d4/
sGLMhRXFHTTGGj4rnI+cioaj4BI9eoN2CGg3O9BbzZKDGnIuCCyiZAt1ivn4dbcV
KxTy2SCC3ugbwPn2AmKqaR3FALT3Mt/KLoznmAK9J25T2AYnI4NwDH1U90e7fHsu
ti9plh8QiS1eLR0HUS8PScqoh1RkvZFaUoe50WbWgEJ6G3ekRDxfha+nNtpWAY8l
cT51b6QOZrpEaTehvqECYaar7V+BSA17Xe5VXwFYHZa3BkFJdVvRNDA1N/BypoT8
KYL/RGEuTWSUYuPdd4IuEeJem6ULvuxmuAQBW7HNtuQtUc+OVnomC1p1Z/T3StXy
Uyqu43+tfKKNIw+SG5Pv0Qbuzb01GR0Ye2ybNk8gZVIzmRwk1nsOG33n2m9W1bMo
dU9++i4QySwTHuwCos5s0xaegQOhtVD+Qj9XCKrwl2n5Q6ZzKi7immUW35lpXWNY
JD6d23f5J4TrcepBkKNPQ5OmfgaTd/Ujre3wBa8SLDgXY8y/f5s/RPx4UQnQi6Jh
mhCDNaC3SUnBDKpW2QTS4W/sdJ/0Y7EU3OKYpG8/ybbz1IUf719fHZY8nih1ShYT
dw62ly1khkSYb8RYAYxbnl0wpbZfiUPUHFS+XJMNbAg/zWOxxeeDGIfSjsvmFFx6
s26sAvRIUUd8BlxjewH9Q2/IrXh6CKFOUt2XUSiS1KIA3xkPuiWL6NtFodRZuRWC
YL1bYauD9yM8St/BYMncOMvH2rWRAqmFUUfJ3rx7letlBUVxCcq3gcm9kVL9ECNS
dKSZivSqlmBYq8biFwBK2Xvz8GXVoypd4F18r26mfjm0TBf90CR/oRBqTww3l/nN
FVp9AvysQ2kPbzqv62dyKGEMpOQM4UyN/iEt3gB/JBp6nC+vA0NcF/i71JHs3/lJ
uxHAAZFgxqMnGDlA5Q7eHcW0EGcwmPr5l2P68rEvBOOasg7bPkiJNvjIJkvL95fj
/4LLNDoUWNd90E/Q3sRFY1cUDEDOV5sgJA0Mkm6kxXFX6TnUelz6u5JgMPHFPdkS
wzljfKIIQJO3eqdTriX4XSaEL+hx9RGIMlWTO9R3sY2+TfG6kFwnRrAfFsHJBo3d
qWIYmMMc5wPuatPDfSIUdCVhcQe0h1kOQyaQ5IrTAfXENQcrh7CjIvhUCIkdXKcu
mTmZSvVMwIcNLIGkIczmX1MvC2qXmlIEwaj/sQErc8YOUIc2uSwiWQEU0cpNn7By
DJl5v9BEigRmftwVPCjXL9s8FQ/6ZQUlDDtcUdh7IYSHyt1rQPul78SDzvT0VyCi
J8I8Tds0If1mD5BdInqN5m5YqRYVBgECPPAtK47hSEjCN0islBE0NkO8Mq/1c/6d
royaAzb0m8zGy3eGdmwbTPLU+mFvFCsUrQZhCyYrW6gtn8EoidkKwmuwCEDPzUSg
NYrzukPDe4bqfZNfGnnKki8Hjv3c9NWvgWz7b0J09oqt8mmlzS/RICmXIWksi4l+
HLkjkhir5SwS7M7sZ1uEBOxB6lp4JwAUfzwUJdi4hfKeysQboXwJ0mgFGEMjmhyB
Ky9zKzTjJTAdmJG+ohsgvkpaKoM0tspJYo/DWfVGtXjA9UttHwS0bZn4X3aitdCQ
QhUduDWdNW0NsKye1c7T3v24HzYPUQyy0jrE/dHKc089SOyYRxXL2vCike9eF4xx
JvUWm2IBvVQHpWhKScxs+XJ5HUtDqWoc2DErYr0lROJVLDH48jwimvRC+9KEtEOD
oROGYAm7jFeGMhrTmc2lWu8O8nVeM4RcME7EGHPD6mbKkRvdgGU2dk0cvthWF7g1
zWqEGumjTW5d0+CSPQ/gf9yEKAuCc3D6NBuJTxXMojfX+Wm8ceng9+zAXMvNpVgs
kQ+5VbDwBVlrH3G82ZpkR0rvUByl8dvineCuaW6CVeAhVmBvCt38YOAWgXvyq0S+
IRM7+3583CMWbnlVRaMYGhHjt5GPBhDCg3nG3XD+//HTWsqnhEOGc2wDzqgpivOm
25jxMeSWmHRcFDUSF0x1Eder4NvA4dYbG9VGHzhdKMmpdvsjFk9+1rNWWDiuGJnJ
2pj+xcnpxckoqZiVpwz3vCObrCToezPFVV19uYstHEOkhci67/8vUSw+RFvEKlf1
26zOd/uhfFolutL6GoY2LnfzT2BvnPMOEVGTao9xSI9DdsQyyXBEuO1JT/jd8q8f
LsvKcESp6GO/5Oe09M/nrUaesbnG5jps1l8W+D4SLgMr+7zWuktMWlZ+ZeyN2wwE
hUex+wUAEKP8ryFHwQLq3wfgP87FujCtqZCJ30IHLE/HAvQdWVC7N1wIV1UrixoK
kJrUk249wr7E5TzW4ZN3wEr0sd+VVF3CGwJRIEoVVzbxsDD+vdY9JbK8xiYEVBsF
7tIkEl2VReUKPAp0+jatzsPs1xP1Kdi72hz157CSmz8gvDVgJx43++6p1TEnHNPz
q8ONyhV0Xu7jLED/TM2uJQAuN/Ol72c8Y6JWis95hyBCQRZ2MBJUd4ISGHMY/5gp
lODofzvhq/o3ePYv2523lpFCPhI6HfOv0ELCjbOjyddrw8THHJcvVf24Ay7vZ5+N
Ca3tCp0i0Z17VDGC0Zfurd01VR2SwWsFljrlaiJX0SkMQ/ee3KLrJpNEZBC87g0z
cwKdWqUH557s6dNSqVl/+lmBSWPglxpM+NZ9K8Z9rS9zh7gbwtER9GTy69WHtQ3i
/2P8hjR5WBYJXGKb6G7PjdJkCZI3OwYGZ3vqKhjVauUKhVPqWP4aRY6E2Y9dW6Ra
fJzR1QRDZHTQh0aVMxZD3yzrsbNJFFcELpuS9mnFQN517aYwo6a0TsRGcMgCUI5G
Zf861vfx1IWg3J3838unzgYl1o3uZUG46Du3ete3PyFKQ6L1uCqr5Ox5dgNAOUYZ
uv+BwF85U+RjV8AcxE2nxQo21AbH8QQfNrxJDmSBuOrTTX40FUNBXaDnFEauqU2P
3qUql7EMKV+fGTgPg3Wc5i4gAFNzh7jFB2ooyZyqLi7AqWPM+NySUjhQTsWFHaOp
JL+U9oXM56hgCfMDEJEVJBmjltwhSuOOJUREYN4vOWvgaPgoymF0cIabJGdjxoNC
kOX2UREpA8/gwbsunMdyQo0V+FtTLEdaxp1RHck7UtKO7Pq2nXUasqzJTzN72n97
Wv8DBZZHuLek1bMgcQ19Yv/8M0LrfZMSevLp8PPT68waqcJAx88qwGRxE8NWm+JB
OPo4143EuN2m6Vkz7GHfXs2bos4xLiYi+i1TggpewLPSSHevdAj0/QQTHbNS3tRI
jrk2pdko460Wbn7M/JRcM9gQhjU7QDwlk6zBYFPmlQ7d2Xst7v9l3JNRowMrHejy
fO8sjZg/C5TyUu7HfuhiNrZJAE7BFWP//vabAVF5pTFT5R3MxutVb3aoBXt976Dp
ImQLbVOw6+vfas29mLGxbvtQNyBxolvszFheSScPTMujwTTKZ9yqjHASLfXApIpx
kGoBHpORsnSdTTlrNLuvdPRqFWOGdyJlgq1nx8egZEGabXWdVwiK8rAIi3niCZQj
3SIqCyz3vA/2V4+HHfpzk2XzpJNq4CCO2hiJNpFEDDQJW9HiEHz5m9DF7OKI8hwr
+6E3ZoQ/YJpUoos0KCOrJukLhMjlMXSPV5Mnc0w/QHwGwb38dh9rPGz20NjT52PM
3y2uYdMNikqh2MpIugHO5IUT2xIEasTW2otAilqrojau5YK+PMvs9oqoqsxuZdSn
TUy9+immNAuYpCK6buYm8ct4smEuEcDSRgl/RUAqdfSgD2QZgu5avoslZhZEnsyx
6znrKjbyaQkmJk3Hg9PzomqOnmkKgx4fbC4za5Pw4BQqpkeIgKWgQ85aD5lr1qcC
tErwAFurfgP3A7ZrV4ru9f/uEXZMyUOEals3j7OUsD4w02b2/vPnVNwm3v3k/dCU
HndIOknW5HzqZHa4Ryv1vOroq/TwKuuRBJ7xPun9zhO+N8IIYet6pPZ0Kjcl3C70
4z1NoKdJC/nqTPXCeeD97kigmpOYkobvCO43uAPsnrQvfoyAmwjvuyzs2vxDdXbp
QI+U0ffgqy3pKVfLK4aqz2B9RRzdTQ1bTEcEmppnizRC+7Wl5kh9rYB+zCCBI6G3
BQGwIVCMip/wg/AfdTi2ucHB6xuIuDgn680QYLwhccAYtqdviU4TWX1wSywgYs5c
tV5iJhtJ1+p/DfbwGdrQzXFKidHKYFjhmOrq4yXQag9HY0Ka4UjYwPjOxFrG40uC
arBMuAqsnJ60V1sWld0vC7n+Si5bu8OkdlETfG7XtRpaKN+WhvZqwWI5C1JyceWu
WVEZYrhABShYgpxb5SlA+Zo2rR57gGT/6IBD+3PNh+7xGLNafEU81JecgI5bHBjj
YJ/Q0pUo4+o9knPgNUuiMK9tcXT7lqgpaYLS3s7kSwS5fVv6cXrWBVJpej/00wZK
BSRBr826lemjJB4w4srlqyRbVr+yUvu9+VL82lAblHNC9I+0/yyaLd6S+Lb24tEW
fHrkWSUsmJUNz2YJisWnB5pMDyWeuVlTXj6av4YE5bP6t9ps6ywakbVnm/rlJjfZ
ZVbVhndqqAkrA98acL0I1DY6ab8VIwzoID0qNhwLoNwP+OtYoGKVSfY/Gr4Nl2js
023d/mM0oooPxK+brmokccHJBeLKXu5RV4etHU4r4+1zNlv+PbNOW9LQHvkRSSjU
Erww9NmdEaWJMUltHNomMLfkrwdav6Ti85lHueStzUF9jAWEpZU5zErLnprtT/du
DxeU8zy4fC8N6xWFGc1z+cBcQb8DOrNhRNKPk0X0h1m2zEkJPH3DIE8/NAqUQnb8
m6Dk2qPvVLnQ9P/kXamx5MhS5J+VPt7x6fC8h9b+FeeMkDFvDSEhHXrAFUBvHJjx
YVFtxqt8ixr+rQQ4aq3k576KDNOuuVyt7HDkN0XV2JiaZvIuPbrSfzjY/W2HCjz3
IR+PJcXH6N8lIgEmb9dUHNNGoHz3S7ENlZeK1N3ve7wEhU5ZpTZFMWcKKfLyZk4F
jonrSrf8r31hupyiftYiQXLw8Sua6j/cXeKpqIsMXAZC+pm+E9ItnJq2Sc6bmhvG
AcV1SEz1h5iYMDHjqQ22eFf8eXj+CHAfhkOqUtdfTixKFFvaJV2K+UUcn4cJu4u+
b6yNhyDpcU9sbCAJWy/w/QNTtyQScNJx0/94y+cimXob1h6l2etn5xonHV6OpXd2
WEaUwNlxCIcb8K/ZU3LO7HJ31grGU/kslLHvfUMdDYse8uGFnYCRL8z16NxHfi5Y
HL7nSfJZf5uoYkiInRa3WyFaRrudgyknuhYAk60SDvmut2qxgZRsdAcaF5395/tD
2iHcudmiQuzW1jJOBcowc/jdZMzWlLnXdSGXJ57xIkIU0Q8V3BsLSGfniPcw/JMw
anQRSQM6vCqvV6NcD6CNRPCnqr/q/JyYXdAoPRKfkMMhYK1HI82S9eqxfmxOskEQ
VhAJeC0JdZkQQd7HnTNqoWcRoYRjpdxo5F0WkNH79nexAl+3Js4vDKz1gIc70gGM
c0jJ5Eii7e2TiviavWfsjVjiLeCVAHqfdFAqD0MzzSPDeZefSL58uw2ZSvmglbSe
4nzcPBIiXdw3iKmIRT/37vjPIJjNRtBMhGf4/TupJbR2bXPSDHE0Ajuvr/om9ust
hvp//1Mi6HXpBNCfJuwvmUfOBas6JOUjuEj79DRChNvxTqYtVwosGsXVO6+9mXfz
hnPZTXKvoF9X/T75T/wzqLeIPGVt32Zm+BBTOGrZWoA5S6MB4kqeKtKGmRsfrJZQ
PEG5LVEy8sFJOHdi6yGXS2CQvMX/P3SoaBdcUbYAMapNrUxis8CEaiQX1TEiUjpp
/QoFZpq4UgbHhKrynnl5UWe2bnpkXap3vfrQqthe28N7kzsmJTuqOd9aP1qDtsRu
bT2pDwcHhOBI+4x4FPAR1AdLUq48PWU/K7l3yGLhwrDM4fe60soz0r2NtA8A0kX5
8uz63OUBQ0wintkeCpcs/ZwLTJt9ncJxWppuFHflA5vnOm33Z1v5fvWbtNyKEk1m
1OvVV9IoEEsWBCSAlm1IsJZG4MfofZF4hradkRrlanROd/c1X+ZYwLnZ3uvd8gmz
YesAnM7YGjcIpxcKWxDL/lKREoGyue4M4QGLiUg2GSy/nPcLnFpxpd4nqewWeuyd
DdGC61F6+ZlW/fdFokoCGW/Dvm0b2N94Y62NGfh75y8/IjMhJoqZ6APPk58i3ZQb
QiNDG5XvJ/oeL9vBBQvoqBqLzNGGgke2iExWBRCQJFOmcKi44XcLGMq9LJSM5MJw
jK4zvE5Rr+9F6vcP+wmEgHCYgoIWkBrvEQv/1CxC1p9Ug28ZGUkCtQhNFcgrs5rB
Ds7ldiHUjhnl5p4NrNqVA77GKaL5upctgQCjYMUYvcVoE/qYRlv9SnaBl+DqCxl2
myie7VpqOR7c3nV7nBYhJQML3tubkR4jiZarxnVeIULTgf+vKvNeNrdwS6rF4ctb
eLh8LioWRHaePzYJsUvpt3PXUzr0FrnN7ASY5Q4wGZ4l8JyblcK+FBZLj80JO1P7
FRuNeCAtqYGte3QTcnHZWg8sLsQj3uOsaySWzGjdVYhS+u3oc2tneY6aqRfuKDfk
xibsFXURZskzlpCrmkmR2+Ql8m4riNLO3J9+aLY3GLc=
`pragma protect end_protected
