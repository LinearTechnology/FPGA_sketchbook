// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ndLTob2OKgF9R1oat4a0XNR4Au5MQT7DezQ42AZKoK377lOwzwi7qKfQ4WYXTKjW
1PkzLvaRdVGpmo4IWAJXtWNli3HBlGeQkB30Gb1A58emomR0Cs+8VvSH+Ofd2fEH
LIOyFAka6E/pzAaZicR8Vd+SVgHg21lPHkTBYe47p1U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57152)
yrSv8dgYkgg+xNGJOYh48dB9bAA0b09NYA3/hQeYj9oZwwAPg81YzpADpN1Yyw9j
SPu+Qxjn/yxigW+MxuS2UIvfRyTBTHUrPus+imdjarw2mW0Ek8i0cPhHV6RucUgL
ZqmtkVG2tr88iV/KJLL2AmIhOCXpq6G4rwSHVfhprQuPLk8XWIHiUZPPUeW21vhN
LUdFPaG9awmLPw1Bb9FJjtw0PpmH/z60c7qpy74G4nzqI7rb12K2aPYrhxN2Nsuf
ZYr64Tnf+SBIzWtwbxWDyxRMDgXRbrd8s4+awO0UmWufxzhrqjkAogWew5oFDum4
eZ/+B1OW5AaFUiVQo6y+B6Nl7zUuaHgjzsgjdQULtSKDU8UzpcTj0JXkruOZekVf
Q0hNjKqMfe2oYhzcE6aHJAxYg1dsYlEYK1epS3I6qRZbYqCBrs886yGecuTjiHGu
8k3yiQKbbClsp9tnHjJ5fFHIzkEGB7Rq1DWwTk7xiDLkTouBEocEW7fy9SWea24Z
ssgjgIM+3wZF2a2qmqNGrD6mVj7ou2l0gz8x1PRv6t3rYe+ZmuIHc1DYhvH5pZH/
xeUStrkxxOYWjbYYyYiGY5AJaytbPvmexs68hRWaPCrLODG+BvmuXphDOugtCTWC
pvYDR67fQSE8gP+vPXTvtFnR0Xhgf1iOuq9F2Vl7rr6kEwycM2cB8sVrdXb80gex
SfgD1PlnsAe+21RpR+Lv6LKcTEl+auQYxE6CvHT6KDgZdOGIKw0AoSoKVClplxs1
A0gNMDr6c8e+5FLo3Nxmffwp8GFtahZdhINpjSgpwlxrG7yKfVZAE8GTMnxNPIE5
68QmFNmMzqAiMp9KfrjgSplUAqePEFljzShNag8BLV52o2vzAizurxn3jwsV5kvq
NQX9Gl+hsxWN3RskC5XK1x2s7DrV1AgdFMwVMY8euf0h80FOsYRpqkvX/Y+R8btj
0j8ePKsvNng6sleubw/6lZRykuxre3ThrESDsFxQxSXCNDxnroLl1uDxQB+4NWQz
a7+l0VPcAEEabWUk7IEHOBHpTRJcP0NsC3GB8UXNFuDuZNku/hKLbdyet29XM7gx
4ZHlfR93SXrE7U/OKmztllwCuJBFaHmRlbotQQWQZFj3lhrVoWtWms5Gw64BBRLY
1buF+iUhJ3R/nEQNXnxQ0+nvsOGjhKkDvdkSZQJl/VTCA6dbGdKBI5bbj6m458N+
Hfkmv4NaBkgV9T4EzW+WQITX87xLEfFZN32cgFTqjDA3d1hDZ0DMsgA/ZQQvtSq4
WL9XG0Ma59pG1p6xiFEAC5LfJJ8b+uGBtAzyk5fcEZCY6THZ6yvv3TH8HaRrTfkm
rKiNxZqoFb+f6zdBkRrGA9ogko07mlHpnc5tjjNxfs33jTv3DeDe7vFBWsiT5puW
yvv5BQHO8bzlzbMIfak4+5GyVz9qT/WDdOFYKYE+cf282PYMOKxIn/6s7Faz9z+b
YEOKO4b30GA/WSw31nP8rztS4fzOqzaEuA1HqcGwDyIyvsqZbPwU/BZ2jcIH8IoF
bw78wkfHBWkyCC5mZp0Wm0FrE1EWn24HcN7phbRXeB2RlN8Z+SbPEZ4l+oYT1B7T
DGdVssHiIwpECwKcHe9pHKFspS/HpYKb8sy3/rhmNE5UnM5phTfx0EpODl3KWuDM
OhHHZQHsL6f7g4ITT9FgLAjBvoDkK0qIOriYOeToLvqOrDsMSGrFAWP90GchbmhL
/IYErFofLdHBYJuAvM7lA/CDsSdVoX8pR5AILQCshAJpaJ3vVwnx1kD1nXVummzb
GBIYMmQEcUn4FxiWfroxiPHOERwLmNNz8ewttlPvuxl313y8TftAwi1zxIzAytPr
nOW7bU1H/LoYule91i86NnXLTWRl2lnhtZUMiQgN12oYOfUSAPD9V5OCQZtdTE5b
JWLhnPLYCqzoqb92/ycrNmRwDU8ZXVXL1RdzD6bbzsQrIv7nz+UO/iXXXl5tOqlY
4BIgl6v/8ViTMAdEHZXQP7lclSQQkQvxNIkLBmDYca21wSp3aFIhsYaLgvQY6yB5
YMsB/UX44VM0wK0qkpW+6Ye3pjJmhTOcTUhowgk8jS+olh7rgfLoWg5C1jdqbmup
+5jgKDQYIQiKE+XmiJ41tNliVdieqmUFnVqdnkcltf6opLkCm8h2SQxPaxIMQLFo
dTefBTEI65RiLUhZUeSlz+40+GHAJU55HPTEY4kNrJkQMrRGKERFg0oKFBbilt+V
3v9YsBx0VFWefZ/X8NPbR0E8u0oIneBZnMOc0VvzikMni9DKu9YfAxgR4oBTHXw9
S4ZIx1j6tf3mJfiiWAU5shNRcdmarjfeG/E7VwatpzRAbAxRLaGb2UIn0eQPeDqj
iPOg4MJK2aibufcdzksfFzKvQPge9FJqGZM0JXezJZ6ccyvjoRoBhTCxWMD9WHc4
IkSPnZDOOE6kwmUQzCNWTBCk8Qkz/bzcuy3yrrHEHy/K41OMJB0Sui7Zq4Jebc8J
1AECswkv+TsEbIogaa6ydoGv9n97X5KYtgTT/5AsFksk3MAReC5Al5svsV7SHvic
K0qMQ8dKU3AMFaO9ApDY5xAtyR0HujZiINEDnd6RGFsP6gpCJY2uVOi44RVa1HcH
LTODczZxde9D4SouJGQYFlz8M1nr3YJQv/42Z4DeqM0psA53gqns8pWZEvp83LEV
zBvC3d4/TGjpCF4t+jhVJJiZObf1v0zQb+2nzQjS/jPmAkEQfeiLZsixSZRTjtQb
1Df2vbmZlMcAlc0KqmIpbK/HrKxaJqLIck85Sm3/XEqONV7R8VNvGHfyMCjduliq
KgZAiPu/UJBbiWNhgqyr6tbuXlM8vsz57TJ1AlZVJPobzJaeaczGAquCkoUbOA6O
3cL0sjxdEgaupBPdfHJuCwsW5zYCrItsXzOoCec6HILQhxsFkPAc0ffxh0NaIE06
T6sgAxDUEOmL/QjweDC6iWA2QbbE//vCgF3PU3b7jshHPn3HXEf1pVimi3qtHXqv
Q3Jim+9yIpHT8Ss/MrYEHWjeiHyErnNJdAOkCkQZP+crcZRomT616FiawVEgpVSJ
b9QBqioRw1Pnzmiebvw3m0TWU/yrt5WXDOov0+tPco7HMybSMzAluHncXjsbL7ql
BpcAfTK3+CWa1uG92uV8oqIFQDBXSSuElHokfWkx4JA1uYrowc0TJL3dpZABfxCQ
CR8206PGHSKrMxpGzHbAIs71qFfIUwXMq/Ad3XRcZijL/Alxd44iLkmYUoJSyJ/+
xf09+hPq/iCl+JighPPgdShL/GiGkIrhdBJwZIfYCLPPe1SHfFuwUB8F+2uo0NvZ
C8OMHT4lq+FN0joaB4pSuFMqVOoc8M7/ZSwhK7bdPv5tdUO1YjP1JDmrvoS7VGPP
Ft7/xTdJ0ot8IrIDtcvXIT03r65TA+8xkPe6bqzfMWMWVvCUaAlQNRChfZBrOTKZ
L2BUxFD5kRHfghLzVqZA0GPxEqCj/ZPKGY5TA7N3oEbFLs34yQRvH2coEs7w3g5Z
V9BeticTv3a0wNJkceP1Xf28TWEdB//CGSfFHu6UrAzGhsBCbEIRZ4yhqeDyb1VU
yhLwr6lHQ+/1ccpqFSF9SjAZ2zySZD6vVnZD9sWNGYQlrVaU2Yp2tOvd1r/w6DgL
JS9jSXz7HEj/dThzP/XMpdl5TMLPcQXcO33hcCMD+juzhQUCTaQLh6JIxdkinGmw
DrnfP62Q/85wqVi7EPdv1qMbl9kdJaXiadJxv62AKNcoE/rO6xKf6hVmsIHh7qYH
dfZ43B3M7ze52ixxNeUrWWZmwCc6owYBsqUA7HWH6uwXN7ZAu/OZCxuX0mHIBpvK
W1wDahiVt+/we3SGIGqkTWgh4FZIbZ/oR14sG50FTeLdutkrOEP10Ruxd+SO1iGB
8Ad1TSbW3I0FzydEoowHHqqVXUMfSUHmIhRDjmkfb5GY3554wv+hBf2353pTda/O
R/rGcsNL5wfON8Vr59o4O1BwShkGmIHN0w0XSpLbjaNHFzvOPvxXsxZio+k1lA9n
8Jzwwvt2ZCCPLghpCrpfn4iYeroMtduO6UXs47sBLxt6vdMNzp3Dgq8uWNHHGMuo
zx1ltpeH073QaMly0FdO9FV4N+ZaJSgB70wVb2ZzOuBYTZcVx13z8yXxgTdCOaFu
Sa0cuE9PIouRjv4+9884NOgq+v4kQM4oJEnNvgzWJ+riojsn403VFm+E5o2CFBL8
j+5PCHj7s0/Or4VhbYi1EAhfGxMdFUkr8X56GvvCS3ypQJyuEzPLwc1v6D+opOsu
cu/kTBMWyUR4o+eNR0gD1qymiXvHNNT7tPIfMkNlxY644aMLuW+HQ0ERWxHktvsq
p+oE92F5/9n6dhRwlJRCdobx5Jp1UwamAPk/jLkTfb/BM1yNXCmO44u6gersJye1
UEa/Vv2o6eDWnaWydzo+zDdchHZiiRQBHi7dOeNq/iJFsGx5FfZp5i90P7m3+yff
eix7qzb5n6R5VCk8eqDdGaRN1zFJG+S+NI8i4xxbopVCN2qWsV3hGwT8V1iozrFL
OXXK/V673vOqTPXN9HYzFp//48gV8AS+8fjsZWl7hgjatZpmG1ImM3oRnFyIQLZh
c3t20XrtVQcy6Ck8cEJd2bqpBz0GKzhrb7xrgXzoNWVNFdFKKkZ5fEwG96HJ1Aac
jSpiK4jhqhu1EHYP2qOmfv+vLKdzv0M3aoxJqJCnRqSbgcf6S7wvbOSrgv5qgy8s
poXjJ3Wtycls/SWQnk7SJrimAl7G6wFnt/0zYuRK56IMcZL7nA4busWQveJ/k0et
ZiRFhl13I56lBHxcvk0BgBPTc3/2yCVoJNGLhfw6Khwh/R+fbU+lxAvpvtTk6mD+
jZycq/OAjN/hG3U+lYLO7AWHWYiwsBOB+jxxgQfw0j3KPLhA6Aqu4gxu5oRcEJnY
J3Vt040rUqhmLR8xfcn1bdBUtfLCNXnKPsYxaTbbBVgKf8BUd6SbW999KhIDHFgZ
Pg7hidPqpQUHKw7gWJdKL1excgv3Fu+o4sJB7MwBI6daUMSh46sT2vdxg+ecTNJT
yEXNVxJ3kBdxlMxWTbYnyfSjV2nGr7wRbg44htPDbtK+b6kEQD+1jLfdfyd/CSAU
+WFx95j1ZcdrLh62BNiSsNzfpXLG1Gi1CSWN/EHf+ZWyIzx5rJm6uS88l/xNhGwY
TjnntPAHmz38d93PLz+kAEisYiUhPuWCMm+02zPhrg2qM3P28OXny7hWCj6cPESF
VbP8N3NlakE2L6H5SttLLZXp1JEWZ4F0C2MHIFnpy3BAFrc4cWL6WO/d0W128qd8
rlDG4ven00ZYRSIrzVsOsK3hDVoBPhuUTTeI6VIoEGaRDOj6LooMfRjQtOwqyGJL
McyMtKahCu6IFCGGkaUuq9cNl3DvHR0S5gh/m3v3u03Ala/9qujyIkWlnKXBWgx2
7ezTWMXx3fxvZGHBuzsYHNn79MOiouUS274iDEM0BX2za0l0MpwJlvIQ9hGS+IzO
c4gqOoJM0ZcWv34Ix2gmNnwcvEKOeUwJhkwcqociRaWNg7CVLSf+q2fBWxJIZC0J
e++A0VWOzZwEykwsx35CrPIeotkr6wBDIm9LvzeazWRdS5gXVQvbMV/lw17sJsj8
jpJNBX4iUYOqjFShcgsKo2iCfY9tSDtAKd6YeR/7YDSPBlna2VyKGyLg8DNi17Wm
0s4uNPEj7tlBvzH6Sq6fs5i1h58Y/C9HVQyonZMg8Yo/mzvwTX386WNsA4H1KiZ4
BGgFzLhakRlWqnQTF5NkK2N+4cxBeuU0aXXzCqOZQny+Nsbd6ovVcr5BDROk6Ke+
vcFXTF/MRLzf6/Oio+4VnzyVk/AsXid4rubMNTdOW5vsqUQXra8M1sMriia1pImo
MyBLTfTyb8Ub/+5RWu4eEAFuhb1yBcfNsRsyiWUKTYLSlCfCjl1FR5WNyzute/pz
dynBbdBkJcvuyKVmNTSNUoGXH83Ecq5PPLZ3gFGRiDdQv0kYUO6LBPe3UD5dLaE3
YFi+MWLC6cfCcybz28fVFq0mbzF77ybT2HoTuD80cK57m09oyMLTFs9jYBN6Q2KX
n6ejSsn3w2wAxLqElWe0nao3/nSV5tqTruHdc8UNha6rr2sQrJIfC9ekItW6sls9
NnDV+Rrz3LV7DWYpMpXCKVjXTRVtF5K9dbMMosKSBsoPhNKZ0cFB6I6JFS2KcGDN
upVS+umoaOMDF7sgq1+o8VNhGdV8C95/W/4eVMXCNA865g6ZSqAPVKaecN0QCPGW
U7TI2kCMSsnlV0fZfAsP53Ugjw4BwiC4I27H4dK/fGmoUPNR62owygXY9dts4nSO
n6R2tCeVsmraAg7LNw308WCqXgWkhS2xL/80cTCulVojwr6t0J7mpMxrRrfv/Ax3
sFvU05iP8XINj4dlPPDwYnK/fhC5wzjAdtCs15vUXODl1HAcm+G/2367oJ7P0qMY
SAnWozuxjhiIymIQZj4Oqoeggfq3Z4mv/js8kBvPnzt34HL5JRex/qIVYZ5JrrU6
DKj40SQilxiUtwt0o9B2NAdvsemsL+hgGaKQChQtZlyLwS6VkPB2bhVePumqiCeh
/3ShL7AvYNxky+FwHJ0DXGaMYwPT4P79QIJS9r9/b7ZMpCpYzJTtv2AnnyhAFUsn
8TcTz/ULEbKnU8vZJh0EccvJPcyfgf17rzZGjROGK7o1CnBZ+mO8ckZ8MC5yziCE
667N2iHEC4UGmjRMRgmgWKSKNrzWCVVDMk5VAC2HTrPp7Lq0CWosbIuexatluOS7
+WvKKHlIq08LEE3q50xHYPS25ffcRZEX17trJQAyq31sxPsqFE5IFu4w+dzsRWWg
9yqdjj4FugkMw6xl98QgdBMjmVAC96jPX7iBOeZ/Bn5GaVZVpTrSNv5lmAmfPCYI
UoaT1e8hPbmW1GMfgMN6gbHiDTcMCWczyImxspR0TCZ9R3Bu8S+fvU19DkoLZg+7
pa+7HTXfSTiZhA+l2ab7msWyHB520vpPKqK+8egVVk3b/wu2uzeIewDrBQxt06/V
Flt/tzH2OxFUU+nGdhcFYY7SWHlt/MNH8YmBixF1V694Poy6ybjaU1C/fOCvAjdl
L8DdItzdwqayNZVlmyxaTof3ryiF6RWuIIiY6uWYqRaiB0tDTU/uMTKb+oEsmsbk
jusCgwGtLNot6/oCO+69GF2ostOW3EDUkiMkksHKO70wLhSGnxIOV/0ozqHWmuyA
JVHIKPNiAeqV6Ui4jLkyigo6qyc9e8JyPMDuGnvLevZM8SF0e/vFNu3oiDbP86X0
uK8XFHBvCTB5+n3lQO3oAw3/G/wrHqYi8ssnatiZ9FDaUjIfCDSr0ZHRTCK/YHZ/
AMMtzEORTs/UR/5o+jt8Mr8hSx+707OYr0KSKEL1zDd+SqDI2qbWhyDgeRaM0DFs
RKmqWFMR23WY0rDFzpp+jfQB7up/55LInTRSljgRQgb0xs2NW7xBCHB8QeqS2tPS
8cl9G4LNBFnOLCH9KG0cycGuWwGVXJTY/RxO50QzfQxoWjZOqvShKLtQ6O65LdCs
8rZNdbsVCQYTM7IYL1FLKsPA8u05OPHCpFp5MhMUoTgX2co9o+LkTtxjm8yo3n69
TeuW7XQ1WvXgp6SYIpndbhfFffVodU8jfvBypagSNiM3BoE1flfzNNArjDBXGlSG
WGBv22webWrVsNe93v/ORiKDj3GoE7nbdNh1lpsa38+5h4hl8ULcJzhh8fQmrX1Y
li999+NI8DmpmNctXm068JZvJT7zpkSUQI233U8vEKFJ10nGUIGez+3tUqQIs6FF
bVCXsflxGOQQ7L3zG1tuMxM8KDQrGmNTZkBqtsw3Vo7o7l2J6Z8IMr1PyCSUg585
8RQegc0smYQ06ynY5elzyNBLlT1LeFn91f5bG+2ursht7nm+mXb7VX4E0T326CXu
B8khoNRCkYVlq2WWCjOviIGpCW5gVgPhXK3XkL7t/4qBS4AZB/jxU5q4lPfNyHMt
O+NCX7NGYSbphoDRpFPTWb9c3+Py2ymTJnHi1/JihD4PGtlYrwQVPfh+RUH64h0r
PBzwr7shNtrMNL22JscQpgAbTN9fBLzrKJVZ8NLy6oSMEtqA3hGdyPQ/b1M74WSx
yww/S0KDy6ZcG55sNaYFOZJDgpX8eEfmZoxxwfXm+qvimVGakiUsajDlDiPlKDYZ
wfgXvqB/p0ITNqpY1Hbscjmnh5CYSB16+ZNFYT5PwUYLPvawxppMXAgjmpqdXy+i
eZsTgMeZyjEEAC9QjNg9xd6Ycwd5w8frUM5uNcISLDLozVyZCNy0+s9LSDliGr8W
fDvoViVtcVszIjnjkkSuJo3iTluugivJcP7FVzIGVWdJ2a3ePZxPQDQHtpceqUmc
mMAkz4dC8vUrtfXMvNNngacxj9c/biEFxEnwTx+S43f8IxydcruQQi4e5AYP7uO8
mVmXQ+LkYm6vNZTPeMBMgfJmyHtm6zKzIMhG+mlPuPkarxrI8Ss9xPwVudo7IKUB
prxUZOziQRjEKOBvs55liJb3o+/kwE6o2KFanZgjxVLDQYTBWX4XIOmY8x5Zodv3
D6SuyU1zEYgqIKwdinHFXILZvAOeQl2QZKFJHkWNJRzSdwzemn8gdE1ZKucMAEg1
Y3qU4Sk36uIksJRjumkhN6Ko5RrcAAAfV4iOGc1DDqan7GVQ2dTu7o7ZVtLcaOBg
WMRkOyLvjqDTsA6W1buo750bdO2VdvTvEmzHsmrVtgA/qupGISdxJkCFWFsvPhK7
b61kHvT4dXBeVqpksoHfxdFYss3g+SKV9DMW1JUoqgEMIwTTY7tpJPMuNIm4mdWG
4yylqJ5MzgPJpvkZg6LPLu01p0CXshvNKL+6FC954nmCIbiT2Ix2WD6Cia9MJtDf
TwiI60Hxoyxhl6PPm6DX4hx4FJEOIz6zwLxWVLcRvo+3DsskKg1i5PMR2IDdHZQP
fL25tRaORoc6gkdo/gKhUI/uqheGZF94ZhBUUdE4nz74oLqfZRYzPijUZF0g8mHl
2PCiuKEQoXNWqD1/3QpILREDRF5B+sr4+IRagoVhe+QI4ngYExG3eZ6V3vgeltHR
X8kd29q0+8TxZJhVzFl/is+YxRrUBwVAVHCVKVphDKCwmxZZhoPfR3Mw7PKRbD5j
04DiDkbnRyirLjOfL0yzK2vVT07lNxD4YgJGx9XgGpTxr4ptGdIe3kkLq8BrDiA1
9JaLfFabVxjxxSvelmdLPjwrPHPNCZ181xb31JqyYucyVaazUzgFBmqkd2E/z5aN
nqyiAbEgvlV5I1aTQiwvbGpbGnAjUKPakvv++83M9WgJtYMFyh3rtnHmYOKQwH7u
AT4RV69Ca/FPY19WuaJaHpNOezJkriab1Ya+P+PQN4ExW+/vj84jqIk3i9XLMrBG
rqUZucZesqfJTFvQzp22eREtP/GY+ozrxXZ1D7DQk5dD7RDB399SLiBSB9lVHNw9
VMV9p8SOvO+jMj+flatsbTi6VJ32scJ1eJKj9IBlwYsFCzCUXVXd1ksxYJ7tHNrb
gKNKY6lzLzV+ImYTBh9c6fDVUCoyHirxT35xKUY8KiiZhDRiwB5kaIeZDIaV+8HK
RVvZzLoHVbTH2LhgHMuInm7dMOnRoYmwcDamlCGHvTFll2OA5ECcp3MF/CzjJcT6
/VLnFAytNH9XFf6OS68yufN3JBzAyGCYDsXbTwJn6dxyMLEONEpV826opkwLbu+t
2KhaAY5NmPXjyrVjw2vO1kG20BEU1HJz+VpGiVLZtYAfoFgzq6e+Ph7FvTx2BanS
YmC4C1yYYSJHOoM3PHAuiY6CuKJ7Zv+GopQMDk3F83Hi3mqHM3fQXZPiBM0C4wrj
t/eajSIa5Utum4X+7FzOXvKW+Q1QSYH2IEIggYcfIDMudgtlGlM2N2f9XaDA8ADQ
TT4VpgB5kpGMKvC0W/Q6O2uD97Hf6OpWKvqB6FWcfADk9ZlXUWyVJnYXX9caCMva
1ollUQetQ72eWwc54MsnfoLGLYGr7YX5C91FSd2kkwhN31UMDya47ymhyy5aasa/
iSbzzMu1VPm37fv28rokGMvo8EPUH8p25tjOiFYB4bh3cjk9JjbkCBA2gK8TokjS
eSWBVNW9dLH04aEbls+f1ixpjY7VtvBYlNmid2Xq5eGsj+sp4Qz0JH0Sf40hC9KC
qv2tjGBC2s1+yU1q3jTa3CrpvdCDesFKStfq76H849Tbq4HXAR/lXBOOwXe3+0UT
oWOALQRd5buFZahwXl0ZprLmI7FVrNySfGyMi92YdUXa0a0iHt8bfK8BGsIiEuRu
e0HDseGepoICe/aZsL+w7qJQf4oepl72ikhRkTYETutqN17tY0ZQ2KK3YISP1nwY
yFbTf7tZ9EunYkbYUC8A6fYxpQAT4ChcStQnsqP270MQRaJ1NR76L+ThxksR6zTS
SCGDSsjd2vJ/LmGmIUXocqdtqE2tbdJ5/QxLk8pqGGdZW1gr2Isn281DgCWj2+Py
o+t2HpXwydo6+OtKRj9WHfA/iarFrLVykiaxGqVkdquXBZkaCHE8J4Mc03fvwfbF
CNn8JbXkrVCaJ0ZU/pvMh1Lx89Ho80kNy4vhpvwYCOSV/8X5sQKUvhE9yyTp5EJ/
G3ID96eMFtmxS0PlGOUYd2cvDa8TnqLpkdmKVKItadt6RlHeJed8qzS59PN8gzMr
upSxHl5G4ST1whBdD3Dsoij25rzqsLcffVDu5Ttz7FjgOddjcRt/liZKPJDNIfHQ
wa5HMtk8YQ1asU8vv8NCAQN0jn4KoODzt06R8GCN+TJsAeNHKvozAGMi7pmYTauC
NLN9RORfxBU2LLm7xp6UB8PrkSsu2xj5SWGuwFRD+Jgqx7CgKy04ZQY7hv8Zwiz8
0vbwOYgEN8oq4Z7DS/rfuF5210BWqlPPx7gKNkaTQdRuFCQdPT8P49VUVTTEgzvV
xoOmvFZ9lXAV2lxpCHKetHyC6Zb1rqN1sMWXhFIm+78/ccf1j+gFLj2XnFwFUZ5+
8b/l/h9Yea7fllcAuEJYJFQpwYlT6DGeHu+3N6Z9wzD6PSQbElRR8Mht2Y2Y0Q8n
/aR8Sd8TbWrW2hiQ92aSzau+3b/JmnO7OAktbZew7ZFhvQWsDDVoesa8L7QKNj3g
GXYrWjDxmDIKg2E4mUDkGN0kF2mT8l9pjx0TlUy1Ge9y2lNHrz2sG7CH3GmPQ9N4
cWNoEkySUXMDqZK97ha8B69JJ3uDoMUcaRUR9sQj7NUvPpsN62Hcp+QMmy4Hk7Ee
F+sIRfNM/mldkVk6YRv3/LauA6xK9lgQNdaxFMUJb2cTa2kQGakFwYu7invNWpG+
SDrDky9mw9dGztaKUQWFdGr+bmr43CUkJMn/JgCNHzAWPQ1t5pixPMaS5xVJGNoo
vKnnSstPTGUpfQXWau1N4Nq92ii/c30Y8iSrHGArgGd4pKVl5nYCJqS5lC/Dyj2X
oUFdmLI9pPMU625kTkcUlaHXIOxHaMliPWLjlOnKsROhynHt+8ENQPcN15ChQkxX
LU8Q1Dbdxh+2//x6li1IHHk2GbSWj54dB8OJhACnUgdBXxw5HPnuOTvdX0eWK4Mo
tXsWaXlLqQpFHCFVjLMmejRSd8Xn2BuHYyRzo/63zXFZGXMgjh8OWRNlVGLA4ynF
TBktvugaVRfpvSjpZtCXj6yRZf6obagklrIx2tL5klGphItRnmc/1GmpL4QqQB+4
BdYYprI8Us7p8owozeLJz4r+xunEB/RQkgeoJ6oUxrMR2+mX0TxuslRoHRaGcCuK
oVsJApY3mTuBrsJYAl55hGfXoDBMkQG7xDTCNNZ3LtUx5SU9B2NsZjHF8y4zDtfI
1hvxfqood1GaAZEy0a7u9cijLB0RYak1U3ULo7qFF8FHQ2glmkwCWzj5DJozOF7e
NQQYXOMPHBtGRkFCld7lTLgmTzcI0HBkxx9b2QYA/nu0le1iu43jbO0J0Z/tbaUL
r+31W3OFoy2pMReZ29jzH8TaBvxs0Pcm5k/JxcaFIsKDSYOBiZnROvltUpKBO6tf
JzVPObsV3KCUqQNSM4ohaz/WQymJHIWar1aJQte2R7rbmjWl4U1Lbzt7SGyDTvUI
38c/TeBJj2myGWacv9vmwQhBUk+4n8LUTCMOkE6OhWYhf/+QIFcSKhYF+uRybSH/
xgDXwVeDUhZFYV0zWFF/axY22S2CS+2hNFJqp3UaYQdbUxR/01JRLYTzSADs6Lps
qgliUbYX/Vgksf2HmxPhcrBfPBPv+WuZ4OTHot6Y97gIAVGuJAb0Afm5fOMFo3ge
8rrhZMqs/tsSJYB9fSgCjJPumE/03sVVlLsjFOSAtwPYh+kgVrWr/nb8UhkwA1J+
7OpTqMZPVsENLFGZzTyEe7hxo+2I1qhYM20wziZY9CxQb6Y8Kx2Yl8VKKzBxLaqG
Euy7cYASX5Q/rRDDwhSiM6zHk2dxEwHXHtD4qZ/msQiRhoOa0pWSFqiW2nuWY1SH
6oYl09bAuPjhX08aQEuYK6nwIq7EFWZDTB3EfaO/8NyKRczXYjY5Z2VMXUs8qQVq
qc3MuBxsxPmHybiq8jrd7V2OFA2hJ/85nSAqhHXtxEL74GTY4gDGgb+Kvhw+Ztwm
pw/N7bO/I+TDDkTX1/HxJzRKs6FXudMvgsY7Btv1U0WpmFbv1N/3u/Kaut08PWqy
SXCTLdBc8zcl7E4dKj+tygVei4qMd7Y7Js5I9rxzcsGbpYE80UyqHBEAR7FeIiJJ
sJYMK3vFU5ldgrs8LZXlQ8CobHXOQ39vH4OwKsHC3xYjnn7V8ktN6tGOWOlR0b/8
O+KiUwCmzypyWp0W6uNmJx9WMgMAGd/MaB4sA5aE5UDOdvEoh4QrJgYSYNyK8h+L
cql40q0/C3orpW4uDdA2gOLDZuTCPcUz5IYlzSTCLhYQjk1VIqgBOO72N+MzocKU
BAqw+vCsg0APgtyTrVpMX1pQ5kajPjswMT7VlE6FXdcofYa6g4kdnQbYvTej283y
CJtZIIJEEtb1DCaC3QPlyzACrl1zVvbEFBodoDH0wHYjfjdKSj+D0hgMrxLDHq7z
NC5t4OwYC0Y1Drc4bAVN84JrF1LUyzn51nmimMtaMyMsqekofTv4BYe+ry43dTfY
zeKZngmqOu5R0GB1h9haq4S3TnSIhJckUFPyhzPcKOXHqM97kfKkBqHyQSBrsW0I
mAPNiEpGhYc8ZK40Y1R95Z5Q28qpJXB24U7f6TJS5HNGF3Iku0h/Ovv/EGSSaBnC
Te+qm7O8Jl5B3rpKKn04DxsfjOp8kKLbrZQ5tSej190vR8CCy8lAZmvSDipCUYK1
UP4APBzEhj20HmQWsBf8BqBFUkLqgXJx0gtz9AOPLB2EWYV8XaxpgXUOeEorSeZL
sq5Sfdf9qChHxvm+1JULIdKXD6Tc8tBqqXR3z+cBK0RoZlfLluhRGCad3Y7X96u4
zTvT+raUYASM9biQpAIeOlmekDVelTlT7wXkxZd4FyrV4/hxt2wPqv7+g5ZL3bwj
yPv6wRxTsMN8hoN+u6XD+ZnkrjHKBhxw6XLjkTPTN1AGHjlJ+xZTAgfQMO5bHsFg
R2Vg3I+qURetdPXrgxA4rMq5Lzn0o4fUAypEjFhE6m26OWaC4LDUxEbcmvLcxK4A
u0Vdr/38FcA2JjfVYc28YzVArT4dg7GCDGM1S8EJKSRBqaRoHUG3dbyRHRdLcyQu
y1834aS/27fYGLGW+/JLEHEVRHG54BGG1vBBVQLxhfulDawN9ZRq/LE48BFee9ZD
7ASnisNYaiRaPJr+Ou1oxIJ5bYjbc2MgrQ24OpVxDfy7uU7ZiAWvtCYtw8/Dvawp
pEzTJ2SiGi3FTSUovQQTsOJCDi0lpkNN7L7CUCoRYYLKhvsxjP5G7IvDDIL28heP
ZDDlEjG0t4wHzBertfJQFD2dkY4tEpneuqY1VcEuTEkhY/vYxCaMoszrpW7PBrAQ
LkYL59gE4EklsgquCg999/jGM7GLE+FH3DGEjFTvvjk8wN4fBIBBbCndfSHv2HWR
dG4Jn2V1k8HfSHi7lCtNHMO50WwevnuF42Tia0p/oThNqznW8TYwolQHJZeygMGq
lBragfdmYtdoRs18r9RJo83BZHxtf1b9X890fJKe9NfIkFdGboYAEXxy6icDlrfF
cAJO1hNAP7XIZ5YZOGcXkDb+ihS0VCAf9HpD16wMeFjiRiEKQ63V+IFwC1JCaiXO
bGRD4CiKCDahOeavn/DwTrncuKOI8j6FEViPBiFwL0Rs+jPxCIdJFcIN61wWVF3b
9M2IyGPatXxanwlwYPWRBr+SvNOC2Wf0MNGpDUtF/gYTs9l+bHTzbd0mKUlE8MSK
hzyTH6vZTVw3lD1YC/JJh3m1mrZENxLAyKp7AF3/aokaQcu1joEhM06Nv4CYUupe
85wukz3WMpkwJE4ChGLi9+f0bpcovxEK7wcvaD6pCqKtgZKnwVSub1CmKbu67m3f
nuNcps4NZ0rbPXA6ceSQGTPGXRQB5O0HvsvF1TAccPAHzJ6RoCBsvOUhQ4K+c6Z4
NEK/PspbwS6qexC7aC9SHBI09muhgiuU1UL+aQ1wYtxSwHpBf/3Zj6UqAtJ38Dvw
dl97nWjzQh/q97bs2tY2+fjZa3RpEWts7tZekA03aJ1xMhwuIV9ojXo6j1mAesq5
n0QuDzrcoJOLnfIJoPWda/1ykIsZntHre0Vnz8APMHAVPxb7SNX3fixqBRKUmg98
eBGa0RUAJlnKRhJPO6JwygAPfm80cVW+5NgKNrZ4JzPtK4i1EV7FReIWO2Tc8Tlq
fX8O+7uL43z4D296bhvME0B7Fj8SpUr63JYoCcvhN+xmagtGlFweVYx8NB4dG0ad
SXVQMGnBNXUR1Uep+Qgd2zfBu+p8EUWjK31H/8f+Z35COmjqQcHc3bQM0Z/doH9r
Ey+ZWB8Mro5qXf2MN8q4a/fmjIy6Kz1iXPYHEfUoT/IbPggdMMrkgCOeoF6iYdyu
gpCmMqYy87J5IbduxU0l9i1Zf8omFaAfeWqKzSAB0+K8aY1T7VIOCVf4HBYMeTI6
19cLg5Mb/4l7e2zfKrbTFmphknwaViCb5m6xOoX+tPoCRzdVzFLdRgyeujIR1hKr
rRX1PK4y6uwGtjVHT2FT534iEfiwi5DCRvCzWxAl0U9p7HgBqug6uWUE+qjyjhP2
yOXQQCZqRlBAdUfBGa70atUp+rNXXfEEpJR/lUVPFADIfX0TF1WEkztN7hMeejWJ
gdEar9RlEkZAV2VG9w9VD0oHxMV+xwFolTgk3cJ31Ei9VvoC0BdnJjp1dZDrzsXI
YMUXSnuFQnckWJjkDz5Ma8K81YWYjjrYe25r0uyCMV38vt0XW00ZC1zQtLLDowar
MuMB64ZN5SeVPUwJ8e8ebCpr3q7m2BtpbYNE7jCY39ZeUzknd+aPD07es9Qlffpc
p85WXdOfb6knXruXB9jJXWXd+kisgvs6XEwB6hen1UfS1ykPmWiRo+IPQ5IMcRW5
GtcylDCvlwD3QRRsbXOncNn1jqjw70MtcU4Opa0rezHJd4fo9E6XRyxu4GFkKCmr
6W8amak0b9/LiUFW/UotpB7nCKwXsPfHZpm9UVmm34yJmjnB8dheYEhsIoDomHwf
oY+mUjrzjWEkv+/VnnWaeUvRM8clSjQ+nQODsTMGSCPhiwGHB7WgKhCs5fmLL1AO
bBhL88cMPyhd6WaMBWfMhZfvyIcm+W2vsCe3uTyiV+BgomWqduSBzx1WO6CUBXs9
9ZwRQkXbxdsa0K5DT9MyK3AAOe7B6IZquQmL79pqEjeyqGQnt2qX+ISGr/3fR2Bw
rKT0wenmCzmNtQjOxjDZb/NuxvuFMD6HmleidwXy6XVTdQ+Z8svkUSRIMzRvDbSy
nfSt6pP/c2JGscpEwx45oCQkG+4Z2BCDdyIl0fCMDaMvSjx+vAxCGkdjad0GnC25
PmIFIqNMac6eqyWmXaIMA+7lj0PEXrU3+DCrvIy+RgW3l0rVNFhTLcLaX+7IdT27
5WpJzh6OXk4oeiRZU5TUWc08KLipmgALopmJoE+Sah/bNvkykUw2IRV9hew4uE+K
mnCL81GJXMExtXyacwQbItg1DHtSw+ZZPgYRVfitOLGOkodWI0bORlsQMsS5FqIZ
ztSw1GTKuCy5OE4YNGbMZbQ/GF/Dmh5ubFzI/8R+tSEjdUJQqZDBpt3jKBBU3uKU
Z/vEAN14SMOYPV7+uokjl14SPeGSxerEWC6W+nAK5+J7d/qv4sA8UcdwQsbjWaMn
+iWsgQCOaEEu/TpEgqS1rFYcncO9UlM1MNDNMDFnn23F+Sa/S4/J/NDz6Ip1tNtD
tnTZFa1OenH5+4Dp3TNpyM4JO4a1QlGI40s9IHRNEYQV8wHXuWbfRHExzUc4dqmd
tJJTRbS8eHftF0rrhCoYddL7JeLZiDsD59k5FdfYFlVO2kNVA8D+wiUpsWjZqus2
+68Z9GGY1z6gQcqomwp2azG9Wf6TN7r4dQbQayoYt5w5AInerE0fJwZULv7DHwxK
OrtzPwiGeIqc2zHVFYN7IkljC877dzh8TjSkhwPIiG6lu+cU1vuZ+evJLyiumf7g
ugN4v5gbxbCy9Td59QRW/uumhvnLw7IlC0/M/2KI9bC1QfYsjzv/2vbYhXVAQSOz
K81nCHSb1tIGEf4L/E81i7Qvt02WX4Vu8QUtrBBWcZ5VJTvVieFL204ssr1zaF6n
kzRMyrsmmFcJEAPnFFoxKq48b7IOEP+FH4AZA/0NenXTZ/ZBhC6sx0Ty6DnlBKjo
pqT1kVOvZWAZoKgIbs7UZpVJvSPr5qIu2eG51tc8oR23FdwiPF3k/jTZTgGQKbrW
Qm9ubXJ1S3s3GQu5y4VXKgQJD07HfppFUyDB9wlvIblaRTYVwrkLMtpKVUUS8ib8
2x+zc7ZwxYuGBoAj6OF+VXnJVsWLqwn0UxQQ1Fu0kV/Yi3zG9Pxf87ITuA8llSEb
wM4LxrutAL+CgoN+QEmLM7WKGqQ4M1NbAkJfh+SSABB7bmfg5n+4ioAnkn6Qi7n0
VkaJWtYOU1VcMF6wkacOdj/PtfpFpWlIx6UWdoNVucK3SGifiBPbOErBAU1DKJ2h
9MNFQ9ZnTJt2kgMKVlYmCrOwlvjUPD+J4Nn/jCLv+i6LPtKneU8uXwur/WdyLfzz
R+XHsRqcpScTWghMBzU2HD7x/IrWxayAU+r8kq071kLWDewUQpGCHUqU0likzqPR
w6Al3igNB4+wa+qbPgIRQdOIJkoq9LzJzeHpzvpUzSVYQn1iy8oX+lQ/ogt9GA0Y
JDHb74pLr/pULYxbHELADvquTR52ttpXqHBHkO8XAvo+fTiaen8G4Sma0XugwhdF
AowLsmSD81Xko8oClurpaERy9iMInBQOnNcaiVDWoHxpCSh3ifxqAbSY1vbk2TNR
x3rnqJLevvbMv7xHugTytw7iqVRd9FhQ5dB/pO1xjlGO1qpfOhcNRG2N5QXukb3+
IBpU6i9UoTksoLLYUvrGGS2vP0jdEs3yR4uxS05YAHPScDvEaePCdy7xu2PGS7XB
fW3lreFr+8w8BwYr/+sntn1rHogLTA187RDwugIjagwJ4LBxNgP3Mnp4McUx0z58
deSz/ky4xBEVLNjxoqtRt6tmhmXq8UxeHC8/393a2Esy5BlSvt0kLIycysb7/g+w
gEeguiB0tbbYlZ9YsOcCRIx2zVKbN6Wrj8+ow/NEPlkpFOErLLx7cqDu6VOEsBDY
UbpKksqMgkbleyxDoNyrgtB0uyz9Ghow11mwsas1D6gNkjGygpNeZdhY/Mal1ZE9
dp5MzXq1uE015nC6TSpMCeIrabepFlWXsh354INSPRmWiHVDcrBOrkW2Sa0lxx4w
BqXBJ56ye/v7RznOSbIoXWcALRnEJ5fCBGCGQOmwxvbadFVjtvc9xO85ZCg51kx9
srfbfUI+wgrPCPDNPpya9NNHPp1Dsf1ceWNeC/c0gK4W7pv7YAihf1zSlC9K7GNR
GE9ha4v+TU1yq0Xj98nKm3yfn46szZyw9mHtN+Xl+PtcjFLnF9h0PdFS+3E0heX5
QzhpWfDsd+DN/43MA4Xy5hiLU5FQ8Ajc6QgIe5NdA/AZIcLjas5pY4QWA3yM7pdE
h00ksEWLEgKHoFf4NM1T32RF8xRySAgAf53/zFsIariBL157fTJG4r8+TMyUX3rg
q/ck/qR+vkh+ZsiitC5c/mQJdc9xobEnHNTOggLwwQ6lZXt76ByCzqLzumSmvwmd
kQdpdIB+L7JfAciTw/oUiKMGTZ8QldPoIRAMaXxkB7D/tBitR+HA4qNAzjydftxW
Et7wNLY12FREQAWdxUh8hx2PxQJhstzwJw2j4S/iUWiVqh4To5GVdk4Fmg1c8INW
W6z1IOV/VRJyrlhCrhmqHdEszV7s2dypv4Uqjsdgot6yuy0Za4WT2KDiDYBbyCo4
p5JF4UXwrKRwLzV2tTx+AeeI31AaAZZhvMMMIDbizfzPKcFUcXXFF4CL2JqGyHfQ
yOrmvsENemWZkPznWII6gw0/K6V5zJt4JwFeyVXJomDC8SERFQd2Eoq9uuyUnIa9
y1Upv4nAM7SXdVRVEsSbXkWmwbNco8Hqc8olMJwByTyjxvGL3MkD2iDK930OPkDy
RbYYYQDrndefvGNaHaBs2nAtS05ttApWEBd+tnvHPUy2+ZW7wHCqm2zROY0/N9V2
C48phK2bVzt3oHYyA9M5LGtctmVajnOdLWJt9Ibd/TR8Z8d/DY6uy2+LBf3qXOxO
WD1F5KItZOjV3qL94uOZWDw2LqPFEkWMqA8BUkxFDA0WMvTrJOppAQUEkME//a5+
MmnYUJgYlBPBtz2B0eia83Qf/Ok5B4xD5KH1dNoeo4MjFa3ia5O+6DyMBkiXtBVo
De81SF063BKoJTPwzG6zB8ETD5sBoqzcZb917+Q75pQZLKF/AiwlbxeBpmQg1/Fk
Xl9oaAt1dyPWpgmd5OUP/rwzjOSRNmburKLsPzN31zX3vj5qkArBh7UQwBHxclSU
v6wsWT/NHIUcaZhc8YMJFSz2AWacEPLopXi8YJTphoU3QMlfwDigu+5QeB4+2en1
0wDHcX7m1IOAi0qfwqsV6MPdXR7okAb5flvFKYJUGE9E4SdUCNrjlNpa5NAK3hft
FFcfZYeFEL0Qwtfku4NNhY6H1/ezRnrMKBDoSnC8J5Loka1KdsLjGlhjRmNecbX7
pz4zIiec7ZbRObmdbvJxiC4olRNTlnq6IiYH05bXx6ndpZTrwEHJzaDoxEOelypH
x5jjxPwILGuLGsM3O2kljbrfw5PKZrx26jjLRdO8jFOo9Su+okCJ3bLePn1wvLy5
3eSeeOwCzcPj8DSE3Nk16HJuzmQukrZHj77EYaQS+7hfSvRY2vyQ23UoNbRjUH1g
Gi7B+rtYAwXL11m1eN86kYTDhXg9no2zVv5Vtbs8oF0A1/fbRT1RtFkQvUxZ4ium
y/8i5Jt/59GPDv4ocdedzqnI+qKO4Bd9ZfFT2kB3gLJ6CZeXwempksEdl7mPeUvQ
drMY12wpHG9xtd4sAs6nt0Qi/thm1uMDzo4RAkeKFipu+JJHgiiiO5838EZyw8Y4
V5PsSesBNPb2rB/A2sFuvMhhiw6TYNPR8UIdyziKte80PAA5DbfcMpENYtY8g0OX
FfKgHKUboQYfjpeb/ah3RuDC4GPKabzIPQqAgz7kXprfDzp0YpWkpixxJDhwbHPe
QMKyFI5n7xO75FkfGsAFBY1BQxZSRGp/l2IElenTohqlJYh1YOrKgTQBVz4969mk
PCWnSw92yc6xp+3p/1L2yut8joGDgvdX5EsaTFuCXhpDhH0eYCBTHaKKNte7yaXL
q09E/nN0BUFTnrZs9A6IryyJswX5pE2/CoR+UmqWwPqLCVfnZAG9fu7As1rAPWlw
ZbcGb4aIJpPH1C/nJMiEORBs+lkjTyQl5NwxXS6R7NSmbazfw5rGCBSS4ywbbwfj
J//93QJnQz4Q2Ba6TcO1tPXPK5TeUYdgr8Yq3Aa935E88NHfQ8qRhbl/rNa6F0um
oB6iU5Rr8WTI95f0bA3LLeo3L6ldE/VmgGr2D071aKsUd/pHnj6+NktNV4LNiBxa
70NB+QVAYWdpFBWizxSfOl/D46HBlCxW58aXUXteHt4K3n6bRxc+lyDEYu7l3hFK
DOK7cnovX//gciF4//yFWZeDQyrnijZhtEmLwwWdYnNC5iSXL0/CHAqXFYzsu/2m
qZqrDz0CNfidtFEmgAPcsaB5e29t8JujTT9qqSClcZYOZXMRzqB/be1zv3TFc9yM
imSvm/vf73osJcg5r8+3AYiJNOeiPpIFhT+h5vYMWNoKi4JjBr4261MqgzlGPl82
EOJsTjTyXNs5E+pL2NjwY6aEUMWEtv0mD18QH2vGcnhGQOVDvIWZATTDU89DRn00
b5zN71zDS5w8znqKuvYqqlrea7ovMrGBwlF9vgLyGYGp1HQ5DHyXnM2kiEzec96n
dkH32EgCHtdxJ6vvWbDKXjJuJKUZlt9T2p3akjgEVxRZtuQ8O2hV04j+Wd1QPCEj
KOT54uRfZq+IJjxJ5X48Z1Vzc60LfVVSbHkmCMuSP3551lWDPgjVexMitqu8FHNH
OIrMp0xSifdZ5kbWR7af3Qv68cPJ4AE6ZQR4YrMctgGikXVDxNhTu9GHEv1DKciV
aPiLOsjWVk3fOYD8W7PWbZ1anufl1OAaRPTy1vzhnbn0osLP9sNgdXQMULKVQ7gj
jkmtV1mFweF/wfDYPAWVdUN470y+lYA36Q5FqAkuKP2KwYF94IkkcwTLfelgU5Cw
GL7yOpJSU6AtF/rOHInQ7Kn+of2iy0BgRyrBHYAbIEnqI0KF0fWbJ1BSsVqegNz8
iZAYTf3V59Xu6CDwLluNHZT9QeygMhMZYfaRcOXiK+LeUY6gIuRADRemiwcJuAbm
sraRIptT8Ti/eUofA1BR8vzNBRrZqo+08PnYFwJWpML5ACGsaVVJbtAflHItQAAJ
yLk1myPDVl3uhitLdHeSgxZAhkgzQXXYjxeC9+O85bOKUQxhM3tBKo7LkV7Cf/um
8IMYIDkKH+JiINiC6wZZEKaxJSj7y3wE9ORQQ8HOofSpkSplNlLtWEGnHYqfEC8N
wsF6fb4uqeICgg/L8HjtlI+UTMuIRLxTd6WgXBbSR4MfODq0drLEcGRNOrw6+eru
io3mYcPO2kIGLSd6lxSRNjA9pV8zEvdQHpUK7ph09x7siGqxI6zVpGS8aIyyvWPX
3gncA9CarjAaajjiq952hkiOpnHZXu6i3dk10QZRlhxiV0OHx7eVm1enHq2PD9t6
jnBK3PsaODHZLE8SpZtA0vMEqruNLM+cJXBHPbrZMJCINbUlgka6UZHHUdIxGYaE
f3GWVwyI3WKqH5SupK9IMgtyI7FoSBchDXbfPhcrTtXk7o0WmXNqdsNC7STvizTi
inLpYlUijQzZfvj5/soUuOd1OPTUx1hk9Qx/FvKl39ojaW92uFqs6aDDfmN6O4zX
OYdYELqPpWkPZY4QwbLDWjJO0pJvTWp52zd2lO1f+6GzXRn2k+Z5q4kvHd4tTps6
NUrxaRs8XkvlpfbCG03Rc7qJoE2LN+3y4uq9Z9D1qshilXQq0WHBBgAiASXLLcaC
an9OcQVwPkN5iBFSebRA7EyUF8b1tu4vS1J9VoiRGHphC4xTzGvim5ZyLSQffmE8
W+c3tgOiRrwtuCfNavHV2wtxjSz/dHNWQtLI4ARW7fEuKAzeD37N3WgKfEhrbdiB
f1/r8yET55zN6HJQEex/huZ6L4PYcIzLrdSi7tLr8SuR8r+c9PYqzO9NDrV+X41u
3oOhWooACJYQ5wAatWLSXv9vgPoUtVEvOQzRHYRitnUH8F1unyU3KqxFfoVZDFyf
yzzsySzrI3o1aDekSUZFsfieNIcay+xHB8rnrwXXo+KwTTLVWEd3ATX8OLX1ZrX6
0mTFiPKk4YwqSpm6rqze314S9kme+lSiSfNpeXu6KJMFwfQ5kKkjzKsZ4T4cb9+g
9htyqqhvizRxAIsUvFx+OEli8NAmc2tQxElEBxzZzsaykw0PmNEpdkPBSyC8TTk5
OpIAjlzMhQw2BhPgROuuBA0GjOvj1AT/q8ytr1/r5JcnUskEvLN8U1TOkSSsXI71
iOzFFOCNplVBtg6orUrvmjwJqvEWY8EsNH+2CIW9cwE9M39hZfmN7CZQrSgQOA87
bU7aPc28erwpO9SZK+lL3T9n+V/pZIPxzpZrSYF6P99Zaw6uzLZpCETjmhCwd6Ua
fHnJyiJcA9qszyDHZahogi4VcCoBfY7riJ+Z4TDfHCrMBfjazlmaiPWL0GpaExHz
vIKg39M6BEYJfj23TA6yQWXJmjGrmWrB1SpDTnB8ugiDdz2wIEJef/0Iel3FwXrV
8IxMv0lBTke+g3pDpcuiOesfC/ld/CxkJyY930PFYGQ/1fPKPJzAZOgbaZOinH/t
ChUbAlSoD6CbinS//TjZ4xP9KEFZfbIgDWCNly2vVZo5YTtdNHiOnPk+ZmbfAeX5
V4uBqiAkWgCyUi5QVRe4SsfZ6qjz8uh0tBTWj2pFJfZhjarTwTMXA9FxBDXqru9r
7xKv9ejgaO53kFSCBmqdRyvZG1hXa5Fnl/mjojmMvB90ay8MZ03/1AbPOI7jEWbs
2MD+dOgHuomQ5xASBskNKM6jOtZXqQWReegL1m+SbDpM3UPrUXJKrY5VYUDAVoU1
sYEO692ZEz4CB/lq0utQurzWtTKXNWONhQcKwEq2StYfOzrtc6wp6pQ9Z6XB8oc3
vSGDBD8DoSk5YPiP+KnnZOPhfXfp78ytVULkOFgj89YBFAfMmKz2H3axsqsjyvEK
PZlLpJY9UAfbqnEVypNGEdHLL2yqunMal7FQH4e2jiwakzKLPsuCRK7558liU/Zg
pNowsuBoJhakNPtzCuYgFxvPGogu0m+L3FvzhIRnYYxOtzVCljfkliZKZGlZOs2i
D2Dg7CitALVizXLfN7BYfj5HxhImdLCvx5GP8g+ChUcnElARXq6dc0C55aN48VgZ
XguJ7VuTCVvvtEwiMhIusE2lkypqQWlUqUKIeafRHPEBmmjxDebLPX8rqPoShlGu
iEmZWfEox9OuBHFqHv9QGepIGzUjd4HCAn0jCzkYDxJHt7XB9kar7jmvojVd16ow
JPYM06GleqbAOJTDSCn0Z+ZWa6xnE1lHq68OJodAFJ65hPrxWRXcM6ixf+PhVNjN
u+PO/kmOuFbZfBVjmJNQP0BJZmEsR8kY8UNMo3hJ1F7Vlke7N6PCNiQsbXOB50B1
/k/RAE2v5Z0jRTHEX2Cjt7vqFKc7vydNCEjpihYAqNJVlbSuDhmuH69fCGniC0wN
zxs90XTn0iDUt9SGDaPTHNaHSWMl0NQiVDUYfibpF776NjfXIPNdAQB00cRG/jqx
+MXmhBYlKZlQkW5nxj8h3BfhdI6IOuqjpDKLy1CJeYn7qhNllhVAEQUSABfYEW6p
GPOR5k4Nk8KMLmy3eL+vlB9ksyZeAPmnoYpi5OKau4hxamQsTSO/jjZ9z2lNT5xk
8XFjtiOn1CCy00hoUE8Df56bmhF2NhLsyySA17Dh/mxdzP9yZK72K97RQrrZJ7Z7
gorzQoRm0hn7GzwnkZEtV4KsM8v9FWXR3PCA+YXpnEOJjggoaDjomRExEW2FkyDO
jqU97qSmxxMwt+wbvRLJ0pqVLAXym0hf7BeONKVQ6wtwlnMoUjB3Ki722KSWwDIF
D0XoWMUmwWd4zRabZJv21MOUofRQK8gpbo7dgHlSJ2J1BBcEbGQFOsh+rNaqQYQ5
/iCfvYARxmwMZng9TEI+gmfKZlslixzKlyylPUcy2VjkbCKVP9zPgovvIXs0TiVI
xsqJhCbMUapXHoPOHwtcwlr7jh6sooYYmSmbpErT7qjG23n+MmkPJlAr+oms+0vJ
VZVKwisGoYWewp416viDvJqGTVXqW03QgV/Ei/TKeZ9Yd9fgxNYveF1pCzQVpH2H
9QWg/TP93edkebSCRPnpxStrntQrYFCuQXUPrwcroHvlgWdSwsKfFGkssR/LUQqW
Ovl0ddMLRXba8j1njMgpbYh4LCOqk7AqVg/OnGJ4IDFAlerGXuOWKu3D7BqOOBAg
Zt80QApqtrJDIweP7Na2YkbPsT1A+WwDoH0jYSBzrKuzitJ3eyPPNlCQcLMcHa1B
HjzFmXypCFDncrHMG/SOk3+q1VKkfBqOS6cDyQn05h/P8wy+001zOzAnLEh5h1mV
ij/lMwwALnOZ8yUetxyzL3Hb+X3DUn5zCfPxO4AnZdg7lBHmdOLp7OmxBY+XZt0X
7MBEogtSViVeZ3JMfIrR7ysWYovuGTzRF4ynjbN20Ion4SxblCQIuItO9UTMjTBD
/IjY7DlBGPeJm36+De60VDKdCGUf4SUrrvW7HAaLqzj1RQgchMerMWZ80Zvy+v3X
XpiQjaeJnBx/xaY59hpaU73aGKqrmJ/ArL3c7o+NrybtJncfMtuOxNOh0EFLc2Ui
6xp1IWNUd4chqFrQTLz1NFAcfM9hiRB5YEvKgrVy+mI5US76bZqn20wT9V7Sj+PR
nmfUSjVsIoZwPivPyqhszeqXUJKVXAQrCWfKiWF6uvg8Kt2eUC4BE9rbNdikwYOg
Ns3ehH5IH2bUYqfm/IM4I1s1ZMkMyAXT68I8gmuECHe8Z1hcShElBDodf/c5R+P3
ihF/VyX//aTG4ZW/rOcA1Kx/uXHf2w+WFf6Gov6xObAdz+xeDKUYGW5pPRMQJ0DL
iLeie4r3XrE1NVWYwt11MHsPjsKQ9/rxnzYvv413ji5vzjVDxpcPuoorUePNGRhT
HwjvQu4clgEupiqZzO/47+i+QMN1BpbEezTWZMYtSxb+uvzKBR0+Tba93/ZsNPzx
KUXKSnBrpABHlEuN1eKrFHA4tscTjIw77PgpkKeHB1s0nj5jJXJHW3F8FXoIdbbK
JwiBlF2nOvPjjF/OXvPp6BX9dDD/hmY8UVFRZshOTJ/EvrfvXbnaYqdkdwziSA11
FlOitQ78sRq0dJv/+1nouCmh6m9dMceWMDnWY41L10NzbfmUfTPGISFlki4QzpZy
g4CVuvDIEov1W6A7tofVK1sYHpLrwbuLB52opIRCzws3C0Q7PoJ6zHfsf7gDX+nU
oSkChnjCLPtBsSxfNF6ZR2kdOWzzpTGS067tnTZUYS80qUfW2HoILXnSio/4nTt0
5nssvSHLUNS9hiZvsVqk+keB5QJPEiqHCb69izSl6KQ5WzUXNnBWFKPPpV5hNoBm
xXn7v50vkvpA3XuLAFhHxXOaK/blgIWTQ6dlnsLsxnhbGogir9TlCiNhGQjlByAi
47RWxUyeltSfINNRipogsqoaCbcXFmkB7SIHlALzLSYppqejKeugga/7Nms9udZp
DFeBBoC9C/VAas6JPNAJ0uUnGpIM/hedbo3M3F11RfWdofSqyjwRRlG1T9daR56T
hLdV9nUEggibhTiph5VwIBiCBJldpGnnM9CR/ZXSc63oos5OUwo+rgkVrXAp3WLd
DY0P8gMzDIfAm8wzaZmZHD1s8Ygd0naTrZCaC30lmlsKN0hmmjQC9vD9w7z4hRmy
HtAmL2ID2ZJiv9r9z297q7R710kc44+VVjCsDCOrodutFyikUtmn2YypKXGERV0t
Kr2RIfFq1vQqV6gDrrJEgzJMyj/yVoNSfceJuJoytyxYb6xbjUNym+RL0YlvweGv
02cj9BDY6uqJiJ6tp4Dx0NktujAIiE5MVj0ZqngFk0PS51aoRFi4U13uKqAi/YwL
IA2qrpJcVK3uic34H/87Cy7vJW+hi3sPXcp+Z7qsWDfnJk0KENXD5nFBzfXJBVgr
f7ed9Noza1Jn4GTVnw1/YRUiAQG+A4EZ/wNcexM7BB6f7WnoZrqwGKZ3t4tZAw7h
dHkUNv2oQhpyiZ+eWDe68IpeNvqAGtEJ6XssRkQPum3vn4KpBTb2p5mMDTd76Gpc
hy9984YpXq+oxNgUVdL6XmJi/QNAXGwJE6BFm/wqrwh8UYo27glma3FQ7Rstl9md
h/UMC82UtDiIpAjX3k3ElDN+jaVmjhfixx7eTknqNifa0rlCdVz+qXA1phct4SBZ
i3hDbN1EanBpwsLY5ZbxDTQa6fXrUcZTvrn/ATk+ip476wj9oq7KDtIqyvCfDH7h
r+mzpMADz3KL595uBqnRNUrOgtM3fu12Efud82t6D2j+nG4M0CCVUhJ9VjrAkyI3
Z33AsnP8Q9nGMBu5ElZOlOKAvBtbvll7af3IYi1jaSMD3+EZm8JOyBV0pR8w97X4
Xi6+Jmyr7VyCKbKx5PgAwECBDhKYfZMKghLi56E7xSfAz5gr8rXr3Xl+2e/+Gey6
KIoxHxqL2YHVhyIldtzxELBcE5joC0fpomtN+7t1GGaAZPQxXHJChV67hHi3k/6x
nE1+jJtyzBxZBdZvTXYZgMbmfjQtRSpio/iV2gTpU7Dd3uhly4jbvOk6oYBGRRjK
XLvSrBiBqfJLvKfeLqgq5i+I0SUqgH3CuaCPhtHEAaSQg/ODUYw+ZBmP/Sci6nnh
qMT2QVoLPrSwH779wIxWI703YgGEe2iHCqR8TtQpBjm67V0Y9Yada101YbsR0CmW
2msZhQ5k3CXcrBCi6VXaYJCwAMo7dP3sxKtAOrPQ9m3j9QSbTNYY1fB1gxenjU6y
G+0FAE3r2FjDtm5vhjvs9uY20+XDDqXN3/vMNbOdF9LluKItW9BF8rzpVRgeZULv
2HpZt9TbTQ1/KO1e+odaweiCwP31DM+SmDTNt8vyH4Xs+XEHkOH0k0EU1JRARg0w
SIvGE8/JhiNRIHLb94procdjZfaC5STq3cxMmORaJ5pj6z2Kb+rH7jXiQSOPFKD2
s1MfsNkyYJqHePKnTOkMkQXzSHg+nW/lPQ9xDZUTmZ6cUnrcs3ZUjnofq91VITqL
zmCugFMDM4es2PbayxrqvXeXjVdzj7MWexEC3yDz2xC35Y5euS01KoxE0hD0LVzL
kTtkr949yRsV54Z5rNmHfE+Djfh9VhuS4pzW1iKhQD1vm8VDA+K7yh9TWdf+PgVq
OZSJfZSOShIYHMUnM6KhtBhGNB/p/Gqt7RPJyChjpwBjie4GpmNzptPVfPf1imdW
yx+sROvwtZEmkXxKW5YQLfgNvwFibyMjfxEM8IfqO/+TW7aW1bZqKbR/bQeikTN0
4SZHktDVVahoUUJCk/ELmLp5ajD2RJd2wHBvuJm+zfq3JBIRkv0HFXasRGiLCERP
qaYSp4QMziGk1XJ/B6ZCCw4JT8lucFBgSAY/1rKK/m/BOfA1QrqwHOvGAP0mrSaI
TAsQQSEXMtjaQHtBj+YX7n4Sx98gCg2zFwCpIay3oxiZ8krXwpY6i5yFl6+Go1xT
Em2VVJMMkrnvvEXoufvhlFGkecnySYM1WRQFTo72SVoROqykoME3ZUizD55aFzQt
znRYXD5kn+9KNeEpTLnpOL5ot4cHfoie07/phDUTJKVJcP8a73/aUY6mPnWUHT1S
9zDjyXJwSZBALnIKe9dn+sXYepD+7YhgbywE24nIQi5GuzDaSqRIJFuyYNkaFK9S
7Wog0+LV1dDO0OAIdSVnDr5neWIubuVDfQNyXWk1ihkiW73ArTnh1LIERzwkBPeB
W2nfVsdEoCCTJesHnY7D8LAg51n5JJmQX/P9WlTG3hA8FBb7qgCfTje5wzuW7k43
LMLWnlgrE7wDEa1XgoTrxjrjbNIYwEsAX2ggT++VnIdiEiooM0fy8RYR6vCQ7kRf
S0NrRRYCBkLSKoBzjJgFMQFKhYywpW0lloSxp/uuvBUO37a9Gjy6ehGpjNBj3+3p
KfnhOZNDyWLWBhU5Wt/YVn7vf1DqMkQomIKHdbnFErk6gNHYNkcbaR1DUO0qMp85
KkQWioLQbIQLOxL9nPyLRyjaM6DY+r0TNFFqu2kf8GEvrw37OAm5+u3/a5yRppIB
BXUYycuMazCbL+BeEgURO30Ph4aaZSFJT+FCsd559Jta/QQeHH2FRFcmHMf4KK+y
Rbep/yNsRUsoHJ550hCnhW+91MtRiOFk8CM7Qg3/NckXNdcuWbJ8tK3v+XLlZvLz
sb/V2K1ESczmqoBobx3/QqlAuP4Z5upE0BBAoebgMmu4tXyrMEZM0OkRGtqgum8i
79aK025fILV6Tb0i7D5T2+vwxJwxfrMnr8DSVtQFAjzQIMKRtx8QQrEh2kQXMnFj
9nNfZEbECWkt2+Ljl4nm8hVU0HHunJF1Erslsg8fGWabrPEyzwaVaZYcqtzEkRFV
od2zkikgzHESPTrn5NCRBN1o7/+xxMSSINCjzHkGa6VPJSp6hHgushCCccZNWobz
Q3ks6/2RvxmnIl6DSmDf4gb3PzdC0mB78Vgx4UqL87mnDvWrajU8flS4n5XsX65/
TOpC7uUKl13gphrl2i7+xYBz3Z8qKa5nw+8lWMkpqj1A34iH+BoWJt6kfuXcRR6g
ASzL01YPvKyj8p0EZOUiOt7ox7KVOMUPWY0q9cclAnz2gHgRdp0OnzlwL7yio4my
emxwaCAnlMD3NAUzsgaFKfn/FxiAGPqZmAJaruxmE2oHxE7dnvK+DLvxSx6Fcdgh
4MAmv6CcgDMiuB3NsmuBkKzL8l0iF5FsCeoptd3lk+DGFjt/JN9al20bYgF+fEA+
PjFDFvC8jgbzGSOBzHNPzLA8nsQMadUJ1DULW1b7v5IGoCMjPICCwAJLPF8H3i5B
ozRfeSEIAqYTwhXAt46hwWDPTWO+gl2BVeV0OD1PG9etNSZROhnkYiKZsZXDQLqR
J7ajSjiYZqBbwiCg6qfw1hMioA3gZ3qX59uRlApb5jk/hycvhx/rA2p1xAw2o/eH
rcxBe1iKTPY68UqjV4oJrjvIan4dFbUsHpw0XIzOrEDQBEBOkNyT0fdyl5kfNVoc
uXg+8pLfwpXO8Nif24eOWS9chALlJ1AYmfZJzQT/l1PhNupkCpTOaIzuBpXUNpgb
cF2hv8aCjQPAtrWjbTAanI8PlMrCJCmX6e/N7MlJ89l4mzuyM3jzmp9I2s6Q0+x9
xG823vUsxqcXpkfeJIV2UsJnKtpQBqGoB/WgrgmHUq3ehnomZgqjkHnF3koAT7id
zWcb50I3hKLChBX29vqPIAfkPkmHdv1O4+juHrJuMWgykBRr1Se3MvH9VTR2ZBgS
erCefHyyGdVV6eGHJbl2/rt171+XI4VKL12Ykcfq0jKbUSP6lRJjRfnVs6lfsIW6
5oRrWLyOE67fbET66WQ/l6S6O6lsKj2BWLPSlSLrdXhYL4uOj6uoEeNxtlJhpxEs
CddWzNSlzuzNkCxhEs9Ah83HO1qvpTjoyH/bfG/NPqnIP7ydXNsIe3yvkeThCObg
AHwubC3auKnGsw6b1PEqmMQa8lD/MFK3mJYuGqKwBjJ7D95rWRCbqGTq0QCS7UTc
DceBCEdigCFlN9VCTsuN4Gn4yqCa+6wVxRPo5BqO46r7EHZXykIaklW3gKkOMWOk
PZEnMMq6sb+r6+CrQU1pFmyDT2vN/7rXDfT0J20BVwE5kjIMjVkuZTyN1aUlVErv
2xpkIkdm7pjz+b4WG8lUINocMWihN03psnH829PZjAhBZ0biaHEE5g6sPaJqqPAv
BOa0ZuYCBpbowybOb4UfX/FwTMpkktwZdiI7HV81mIYk3XHNlhmazLy5Jxt5q1wS
YabQ7zXnAVuG1bmBdvYfh7yupw+tg39NMZC/p195mCi5sbXbKIvK3uoC47Ebw7L7
qlPuU53gXcK9aIfj3CGUjgXMyP90xFjBQqtPmdQHMy15Oh2DQ3fwBQEkI+CVVGY9
A39mf2pAI0Ti3FutbC11n1j3T1O5IEtatMkmh3Jg/dMr9bYNTDRfcb7gGqYmyz13
VjBD+fsIwp7XPjBeCkR590D+hinFG5mI4PxJfUigXpZqCVh8HvAOhcsTKoF4IfVY
UYLhptgFFop4P7YcirQ5yl7EBNjXA+ekA0U2hBjdN8mMWPFRpLa4bv78LDJUmmcz
saAUNFeVpEEOU2X26XZPD3O8QUl49z70I27yGbkTU/+IQhen82HF+hHd9wK/8cWF
8Gs1rc//TbSwKjXNcrtJX4Cu4RPuijoK538OuDrzCdGemSZ6w1D5d0RylkAi9mx7
1BsvBHDT0oIh2jDVgyV0SrKzxl/7tzdotS74JYGdu5TA5iHKE0df68E69i4X7lvR
Bvj/iMBz4wm3ooAbcTY8jH5gY6SXQ5UFDMENK2gtAh68WWOzvEzGSL+wfVggf2Wr
aJBr0Q1jhUniIblTW+5f7QNmSqkQKHh5rCd/gJV4pYOYCnjypx2J78g2cR559baO
UAcgQ87b4bNRpQjk0wg3pScqqdd9yLpxQ8XE/gkjpuMpsY25bISbrBvU7+bDCadr
k3bITocVGbsU2wAOKLjWAInB7V3sWIzSQCnILwgCxemYFE4Dp/Ta+yKisVxu2QOA
1b4wF3IjpXudD0Mkfpw4FMszhuyxOVPNGebuZ/e/jWtO05X+waQwgDefKjJZ7P3N
wRw52qc8ytm8G7bk/29kvDwQiYpoYN488ZQFsJHvn5PIUJOwFrYuvASpsBvPKm1N
9gTeOh4RsafwNDpNknp/SEqPfjdvIiPjG2LLmvcOLRJiEERbliEy33clHg/P0OUi
5wGAnGD1QQS844JPogcZdGkoZZN05SUn1gLuhPOBCkZ9QJ0QuTluKQnhaZEH1BAq
ACxz6GEDcdD31s4g24kR2oW1Go5EllumPmR73pVyIB004peeq3coTp4JdKwpPwx0
gDEY7U61wlRuEVu5/F84RFRUZa+5D+AOKg4tGrMucdN2DefmNH1/sqHPTroThdYV
tSKPvLPmlPHy61FGdforbgq+7kHpfRyCoaOqtdFJGXHSOLBjzFdnV6uK16vV8Too
WpWpnIzjabR+n+Ry30op5TNyxVZJ3g7AFSR+NA8+vruOotXwnqpF6aP8XOEwR7Ym
VRsemEw0T/CTR25K7/sLP1nA+qfhMAHbzHvhmFTto1PsXhLvSn7oLPSNH3jVy8MY
KSyUI9U1kyQwsh8PJ/j4PUQ7rOjwKXzLidtg1xVx/98ByqyrBdmPXJn4gxM2Owbw
AS3BUN+Q2SWYk66jaUz0V3A6SRom1wzTgmLp09odmUSPr6x9CMxYm0m7rlInZzi0
InbUmZhNJ30UIzExAMNDUQZL6enugb5PIBMasCPc40TkJH+Q7K9OXW0G0qM64jeI
0Iru3MYf1m5FCWYqAjMhSVHmCugnK57YfYuLCvLMyTYlSBq+vsejGcSyNvcKuOzV
t3EjksGFeMLwjano0rlhZDVJ09IKKh2Wv9OkU3RpAOY500jbj6Tv1dbmBQe8bXdD
nt4N1/9oVwljCCY52FwedjjhBV03N6QajqeViVvO7te4L8F8HOu5LWAluOm1RVn0
LFk6CXy74it7ig2cMeJ6ioSOkvLm1yzJBjZdoprDmymBp4Bsk+lpXFPVhNOg6AGS
lCiP0j++rP1IszfgGl6vnpgaaki0AIDofLyBpfYyKRHGpSUMnsUwzOvDIsZH2k+O
bl0zpFrktRsLFx8H78iM+b3f94mGGIy//U3G9RtO1nAeV3+wpWjgyCgH46pPyfH7
LWpLQGecA8mVMPpqHI7PGJTDYBZZN1zswu++4brm+op0LWb7PvQEvBeu9qYQXNuW
X/EJXi3sqYd3ARfAL5Mw67TIRxm0pzPkvXJOuwJsWoPheBSYIbBxTSsRrFVzHoYG
geBKIK89wP7jGLO995qq/fG3IuSmtepcvecY1S4WxQPDR0UClfAnY2YxyzWbQ0vm
twXtXkm6vEBIqPYx3mn1AnKC3StHBXE/owavOn3zX0eIIC7pbCbOFrhsfUiwN/X4
LBd6SEIvMvguLkQ+n0EEA8Utnp2fLZI2hTiWOdfa0031U86SafdTHfn6QXADnGhe
5n2QzQY47MQYHTJz/2Uv3booFclFVceLHLQHP1hnyrFq6Rt8dD3/gw6OaL0QWMg6
22WMwNVQWXCRl3GRkoS44l4DjUqcYd1lfWBFZb7BD1JWKEb2xgP7wrPta1kP7WFy
lH1KboGCXvkUI6BVLGnYR1y9ujeM+vq4lPHbt54mcR8kRILKQZFSEmzniZDLyBci
U6EW/s4VdzqY3qB9+flhegxCMsAV1FGiPm9+SqwGpYZ2Bd6S7IQbXw96/MgZphPP
Xo+zSUGsv5ugdMCwYuS7YCRVPq3OACX+Z4yT9oDLB5V/J+JdBQPu3LpdFbgGcmsT
MIcuaCsWBGsSMKLLwvVctghADmYWNKrNiy4S6S2EXYQIyzSAGKd331UIlbpEKgPt
plNb4qVX13XZUkhzbdXBCqfOwZzdE/F/0WxOzJ/OIS3uVSqA8HlHlVv45FcmS43W
ukKBCDUwi67wIJxsE4Mj8O16C+1cGXL1FKaFEIgPAU54sbxuOfahQ2pONZciA4FK
LZvwo9QNxoIIe443VmAhHdPYWLkZAEJe63io8+ITZzd0fQwi0L7hiOQyn//GGdpa
pPr4qMeZNvfoD0QWU9iTqMWRyqttaDj/Zcib+33l4gknv8/ZmdPL4L+Uhwf67kxR
+FZpS9LuTkjxdOQZrUcSLxRU6DnL4CvBpN31MjDITdgaPpGQzwNtWIDpeUVWmJLW
wbeZpN3tcaq0dXWRhpM8UkMaj8McjBPBIMerZqGNLkOkS45PxTpDYpa8FjT4r+i4
Wryju8m1eof4+m67dNuHvdzs5jghkUe4NeRzVHqTmefXH78o/dLkhGgaTVcVLNfr
7WCjeWRZPBf40/rro1b27kn+csRUCAJc6BdvC4bcxMSav9pPwlZfgEySdwlHKrct
v4sN9f26peomsMEAEZDo2sq+eCz7P7IiaAgDZY1HTEkJ1XNRwwyjLdncOWBfn7De
ybBDtFCY5ka4iEd/aJYI8JlnQRcPw1iWuifMjb5vx+mcH6Flt/6awxzHxHsfn6I9
pdJLFcxLupRrhGiUhEQOee7/jLFy9i4rRWifyruJj51ndGke3DqDQzseJNQdaU3v
odIdPsLfoMIS/xMFBhlLur902HpbQTSnSkRm6kOCdqA6PJnIJn4g4vtU0E8Cu6/x
zdKvk28EDS0qXNg9YzVNEDXcL3yt8VOa6OC0HlqBBkmP2kJiDBqVqQ1kLSF5tLA2
Hb5jnvI1e6x3TSBKjS1fnk8DfItMY0W9OsA/ZUxGAIYWuKYciONsFAVvrw4vThyo
ptgwuJbDnT4eAd4yu+lpr8XTm0DR9p6jU8ePsWVuxGEnQFIOlHysjT9gKdXVFTXd
UrErmJ1CHL8IBGv/3QztIWrpaMS/16Qsj7nfJdsodY3cb9e8OMQRnfarMlOdOw1v
FOEs+LvtSRwBMGMPSlT0aQB6nyoEi3OLtB1rgaJib0LeVJ28x3Whx01ayIHa8ztL
9G86vY+FSEGFi8jZy5TXGLTjv2BtBqlu6hhynbgiAzEkdAlvOUAHSfx5Nor0q7qU
tIukeFoAiurJVsCrvBcXkzJwshtgs3vPrRrVaGGeoBtiS10qeCpgq3nJ8sJbDdjl
A7iiHobGbnm6t7QVqJhkV7I7AhmkzydlIMQKTYFWWbqq6TtG7j66/UErr8Dvww7I
t/Izc/TwEORkouWbxmt2NhvI3SOmy0Y1FZG9NWE5AfBVSzGr3D8tYFRQgFJI/Fu9
xFWKsYRRRGiAVKvMWQP5K7ZYUAWiaPHACeXe00SKKSFv5SfcpfYFWO/X+8EBb6QJ
K8qwl5WcRXxT76cnuBAlndT/Ew2Iyq6GYDAkX1KZ2FW7a1BAmo4TvWR7SAzEZKA5
glbbZKVsiOvAEU2s4HJdd134nUQgYCO/vZhC6bkViTGbgT8ohyzodYV8I/n8RSB0
XJc1pA/IvOf7PS/AWDSa2EkQd+stG5N3QE0v18W5IU5qEaSXx7Ne/rPXKuh7G7cj
8ODuRVh5v31bhQ3ffA6Yb17YgSmoONCsO38ZPxp4dIsVCoYHysk1d7h7U9ajTodu
lLjvfcylbGpMQp9IGmFXyCK4uI7GBT1VurBvIMAaS5cMpWMxQIwQDHLr/EUrR4dv
lZbMBh9HJopTaqkJ04mv7JMxZ0LNrcvf7vqXNql5KFynjxhrKl3nEIK6fICUS/gi
zDAhl/914ZHmFLyyRY5q9xPvjlPMSVgoPK7yhtu4KAeAzqrmdNu4HiFv6pXvzphx
KUhdp+4hdq+0krIr58yj4mevpUxKRIaKbDeLcpAvwLFOcEzoJAuI4sS4P7OB82eW
GcYFocqb90rA/ygy2f1TH7vx0KJUAkrdRr5CmhDa29zRLNjIvtRa1QhvWGg+7fRK
6/fwvoVgG5wzZBRg2LPbCbr47RII1i4v0UhAGezeDs1Nq/JhYBtKzmpoUe7dUHbQ
zz/QGK4Cwv7mxy/L8GvRFeLi8DzQ84oVFis5PIjcuKM+oMKtWZXMMzU/YN9LU1qT
QU1KyhpnujYPBmkNP7Mzy+nBsPaGyzZ/UaYtzbghO8HoqMei92jzR9i2cPbS2trl
dp5lH9M5UvTn54CY3am9MYAsMBULYTWmQcE9mdmTTiARnlCaKXxgFd8ohmGcoFEP
hpxLwaU0c5Jx3bMTrrIW3zMgI38ThdmxowTAZeqxBsJnAeXH2sjzmwsqCyxjiAdg
JPCDA6NzfcHAmhMsSur10HDf+e3j5Yj4U7jGZ1fCfGIITpBvc44rI3m/PyWNSl/q
Ckj3Nq/gPlt4sg8Ki8LlMmqWfbWCPGXcmb8N4xLxFrut/qgmbUGxSD/fiQO+77ep
zIgSBMVO8jNx+WuPhNVwR4tpzwiNb1W8FBNn/w79lRYODutmFMr3u97QEvVHZ00N
2ixDyIel9uAfDs8T4x3CMbxiIdC5rQOm074HpzkrmmV2UFt6Yvudo5DJ3EG05r1m
ASCZ6haqDZP/QOGe5SrZBH6hQYFUDEf1otylK15xR/NRUCuo6uI9MEkhmlJyT2TJ
bUm09Y6osKZS1p79jMeWuisv8TQ83JCQsjbe75T5TYHmWh2n+fR0JIFbEIerk0ST
vgiq4dE6Mi3VeL2BbaDeZrFOFitVD4coq56eHXZ7VRHW85pi2CE3faENNwjyDT5Z
IKXG+kLJHIwNeKSMk1S6mwgPlTswPw4AOQXZ0F9H5Jh+1IBbjALBtScx24qxXx+B
EhO67HMVa/a6EmYDIAmIIemYfjZPg8iHJzWeZF1QAxkrYQP1LtEv+kCzXHYpaJoJ
NWch+Ii7dwECDvd+y0SAA4ZNf1m+P/2ibcj9IEgboB8oliOz9G75sugi7sY6LMIg
zwcQ2+M5FeyP6GNabsQ+t+l+UoXf/E4QVyfrn4vQG4H3W+haGYSt2LJIR4GLmMXM
7vEtIkmNjCSiRrYOwnzkdD8IM00agabwhO47UdJeowM96SWdpwrXRNmotlVluGIT
ey+PpQasH5eIcENQdno6UqT6KISud7xWsoEbIrZh2PH6e1eSs8XPXK8QpR7dGyJF
PJUqBnUOTwnqV9jc9mIbXp8lgDsvPDt9xSvWUrLqHGdrM6iumXN1eRO7o4ZzEDyN
lTxgZd+34RPEV/DLMxxZOhsZ6AaaiEh44opV3b26b3iNZevhrR6GcCxoVNCrpjpG
5kiiVQRgMHfzv1gJO2oN6kltXD0Qk8IFFEes1ktUFAFeoYaun/icM8FvksOuhiSW
9yknYBIS6qkFrcYd1jpX6SxCeaGFmpUZjQn3SdYjlKIA5pHD2ggVsvZuTpy0GS+u
z1VYgOoGoMAOTF0/wByVPvpOspSABvN43+13owgQESSxLheQ5nmUC9Hmx4j5DtRY
cUDOVWPPoNx85j8RP/QuRdIt2NL14v46znPiGBQ7MESA4ZZjA7UaqeI67CadgJF9
xXjFPD3QrbFWahHn3Yp7MxpoW5tOwbjL5MeIRCfeIGWzUUJBca4KXHAz1JLjUtf9
CXaBSvgCvV8iTNt70HkjgmMwqpwgqdCon0MSOf/2MKeH+pickg686OhgTzfHlQBl
r26LAmdNwF6gwBSGkxlIF05lR9rGnZd0g19i55WysolJvIZFLURX49aVDpH4vW/3
ZhP25rpBAuHoaM8V3/EaNja61nBIJZmIKktHNhzDVw9UMe8TWiDi+/VjIpsoh9Jo
Cn6K2Rr1CwoHRoF8ag86qs0X5NfwrfmDSuV8+S+S3CLFKPMr/dSMGlHLy0/lor3j
iQetKyt+Cni+b+m47/LeszGO4Asaiv/FqedyvZ9e21jdmkx8bMa2tojZd5iPkzrr
npFS5f9wtTAXRJGL7so89YICXEFZn2oNm8OiC69C9Dw592dzkVbJVI6yPr4rPS5M
DJ1s4AECNQdjE8DWOGcauFXC0l4s22AAVAsZGSFQNZyGC1qZ4lHybHT2TIeIWuWV
g3F1zEnX08zXdMveMwYeAqpAVcAWPb1k6Ig6HeA2Y2kda3CM6WGP5a46bXQr2rr3
LFh069TMaypHVmcy3uO+CDJouLw50D3gyQsE0nF7uBG8JE2Y6goBqoDwQEVTqOCO
8dJlZ4dM1Woy5bAjYICopd9NTb5bpXD22r/fwZ5voWwAH2f2JLJAHsgS5R+PVnK9
NLWgPPPu+jpDRaNE3IlVKia3rsGnXPDHr8Jl3LZA+je6jVEWI1aLZUifTSROOquG
f4D6iiwbm14CYJHKrTCXNRq1el/TI3TbYqz51N4eOK4Qk9D4l7rQq3sqMpMRZ7zi
soJ8Qs8nHFtzB81ac3DIrzDhmhRJsZ5wj4A9r+miWPmtfRnyb+i7r23SOPDW7BiR
A3Lro5jloBuEyyYVvRjZkOABxB6WS9oFjQzg4NCE6UsKltkMjpwHHA8U0DPZRU1d
7KoW4BPJG98DyOJ3CJxzbGyi8MlFSEBwWEr/Ga9+LfsQbSauhA2FbniaC+xBQDf6
l6HIPNCesCCCYX9kyiEauLiEOOQR9qmTmrXgGkDNYXxvd0mjDWXT4xjfLK0wm6N0
yR07nLLkAi1iyx59tcdhHSVO/rubm8MfII8WPspNY1XWpNdgVA6ZJJO2KLGZis2g
PuHAhLkI2BGcl3yxXVey7vHuoApXUhhOU9EwoGUAWlh2z+mmPlNAQ2i2pu5OgJRi
I5Thd7DA7owQeMUhxW9rhMo98AcwxTr4mrOrautfzlQK7vyRIvYDwG+LU+TTslcs
tA3dOCAgs58xNmkUnYdQBfxsI0+eekgf4SR/EpBf8r6QLjKZFEvrsOXLZ1tx2rii
9XyDU7nuQuHP7k/BSw/PHHwymilG5dXhrjtBlldriyPK3mX1g7yCEMjOenhKmaMo
SZ5CVwBXyV6ixeWm5bCJO25dsfCJrhamkDyiG8h6v7PUD9y6NvGLiSwTiOAtJE8b
i2h/2UdArUIBnURe5fjoXR7oCMm3qoM16FO7RPDAnZe+l2xaqSco5ycIQckwhX7L
5Ogv6HuBNt1LXZInb4pDL4cGZ9vjU8Yn1/QVElWffwfEBKgrLwKdAMRa8+0GsZJX
2bklhLGfRiUmVsLH7NGKEPoSlW7eDjSWWyBkjiuUOffWaRBDDLWiBS3HZ6uXf+ng
Mw1hnoRzacPKzx0OKk0xKS4iPedC+MVMNHqVJ7R3CDOGUC4dE5lFC28ZaYshn47h
qOrAqq0jC10+fW8dD/3u4rzaj2q8SCsz9JiW+NUvDKfDugNqB7sNvXLDMNy+snW/
FvBVU7JCErE3vqmHe+OXXh0g4RKcld3ow2eWTLWgOYv5zo4VoB87RU3732zhWUhu
PbNCwdjFOKMK0+Hdsfk5fChxo3gl8JKe1l0lZkBLJhVrBosjTwloHymk8pgt5YZz
GhgL249Cmro5PxxGUr8aCnQ7c/6Pria9g++s6ejJEp6YocOB2tNv2URMz5rjA8k4
lDhBTBZv+TDNYLOyUnw2GDHaZnOBbVMg/tShBezhd279FjoQDGUDzQatyC8WkJnX
f7bmaeBhgjTMXC1mfWHfEEqILicBmCi4TTsvsUiF0EdpIQKsCaim0YiiqCgVeZsp
E9R4zZ9UKxmv8rRxlkWFfWyjWLs2MFHq37gboNnPqbZ/ehuGcjIuJeBw6ARzLp6Q
e1oH5MxcwdnRjA67ZMXZZMh9zSrgcYJ9jt/ATnBH/Tg5o543uB67ZV7zrpgV1E0Q
vr1fd5jBgZgzfdRQIqbfVYaN0B4EaQbBsepP1XPWZsPQ6VykKv/3YQwtbLKS8QQh
/0jTpmW5lDVnTqQArKf6A/GFLJ90POMwsiWnkXJrXAzG4akD0uTn5iBEgEDSIRXS
dpEH2g78U1+fvWsij8MexGPFeIRgsQm6sQRANf+sSLxhdOmqHGsWuyTJ+B34hHes
D8WT56fb0HtAvWCk9+sa8aUxLh+AeDLt5TpN8j/71AG2DMioBqZmUCkF7+HpM5P3
HSqK321dE+i3B2Zwq7zqStSPgEHWyFH8yFgxP90Up6zufZh4rdSDbMH5RaoQ+wKk
JDmceYuerayrW89CrB9VKxr4UTGk1QXUu/4iGYf7PZxjFen4Odjkw/2D4WQcanIP
BoabLjaXWv1DMfJpqWtQEkc5Diiklx4HG9t5N17s7g/c7o1hh/38aItRou9PYKVF
OV99WPR/AMSyrQAmn0qxlZDnIN0/hevQJlMmN0IXamYCsFkV6mUFIA9NjB4ud1bc
83X0bz1slKF60HJTz+0d+ZPVbgZkhb+RUocm1qpVm7hT+zsXXllk5f8zv7I09Gke
5Pnjk59UDMZ505vHBisRWxS+Ue1qw3n3q1NHW4w27ZEDkf1XeH69Z+KFgdhLBZEo
GtMDQr+oF/rfCRAorLo+Flaqz7do/tgzsX21EVoazsn5wFVtIVzMp3zgBrFh7RSy
6I6Ay06oAHJfhwgaaSgs4Cwrpv78GjGgdIrf8e/UgghsY6K7YbFns1w//COg41vm
iOwSjYCTEA1Rk6PEgavTLhZq7Fw+ZTVu2QnBszds/YAvFYIt558Nn3aenp24PrIL
SRZxYC1pKY6UC0nQASKR7z/Q6imb+IcREyC2Muv+zqQBRYY7eK43nYJYdN7WHPzO
BUpGpoBGxNGV8fmohnZItUY1SBtIr3dpmrCRQVOoMk+z2NAxWlYLGxv+oRIaimv3
jDdFsDt9a4CLwkbJ11+vn3RaKBoeGaJcwG3cOy/xM7MZ1XC9+oMmzhkrqsEtHFnj
2XYqn+FF64KHnyn0UHZUIqgzbMW7P/DoO1MB9KlFytL8Pz2cdY6IyDa5XZsWYTkt
UG2Ws6QQjTnNGhF9Rx0B5zMOTxy+/QiWpANnjHdtNfaqDowRUs8QHI4i4z1Ciqjg
qnkhOOKSZUwCaTehuqG90twZJIz8Liq5Zaq2z/7SBXT0Mfxv4g6jB8w6A/DZCzym
xRAOFoQUJl5092KlcfCAVlwnKdlZGBnV8xBXyrF/9b+5gBbaSaIN+E/XTExqEjZm
DzWihJD5+cbi2Vr8z3qBEHa4vZHNraXLrX8dHsm1lSJfczUPW51LxwMLIFVB+Z00
3yinHjGTFgqX/I/kZNaRqP2AvbdPMk5Bgg7epF4D4dfhxz1aSx7dF2dT2t+Vhs5y
TGxjMGyX0BcgFwFd8wiiW399ipKdAVSysfIyOVUVJUTreOP1B8zdM1fOjDFgZjdt
M7KTUOaQH/sNXATgXlzFHUDNZiZPxOOcN6RhPwsxxwz5CT841qy1ceamahDlTI8+
MmVQAQ1uVQ/SxAZjXrMbSLDTCZTH+Q1hbtuZZGSxXd6K8WOy7IRElWFeHOnyxPwZ
j+BgUhKu9SZ84Hl43KKQh0PCKwHsfTuNu5a8eQVn6KnQd6rBVg8pAsF+TYrRrYI0
zZ9NkdSh+wiIXIS+FoGYVSWGbsD5NAc8ufjwCwdor87g0v8ziVXQRcugiRSMNble
Nj/cT6FWn0jQusEFZUtuXcLNWjs9iqizxZDyMgUJqr18WZQWCna9asZWLr644/Yw
4Zirn7cBv1dE1ILYcSpNl0z/dvFUI0RbJ1BnBkQrgibESV7hrSv/UXl+TEL5w65M
t5zhLvVv74+xyCewDwIDth5exj55IXi0bRKuxl9YVRofj9EMjntNj1npk2ili0ke
WbxrggD8Iqh5CmlWDxO0CbXzdUJbAoMrXyUmR90VIblXMWc5xtruP9LYfq5vIkGe
U5TDtD6AvRArpmWZUnH7uS/wVqI2k7rWhOdH7cmas29EwdqY7gD+Yz7OfDxaRn/q
fJB5GsothYMpEXzdeaurmuM5mU68kDaNqabAXhJPTgg+AH/p98JuRDkxOTE4TVQU
0ZJqpisei62jS78/8v+ge4I0E6Qo84TSBzhXQbw1cgDGOTugb/8xlpmD0MD2NTtt
5373HW6/BrNiL/P+8UpbpiBj3ql04u9RMEYhh1xelvyIyL7Jy35bkGMPpbpbLfKM
cC4ZdVWF+LqKRaZeFS+ldN0v9cdQlABBOikalcQj8fXhPpvdotuO2SQeNb9Lpp35
Pw9UPF90AGJWE4T6YFVP31LTRFLLHu7w5pPWKXR+UUYPoeYqMMGZKxhTskuo3n3u
ipOzsZXjWCi1J47ENzqJPM7sYrg3JFR3TIniIkfi+CGgMQUckkNNr4r5f5bXy2ZB
mm5OjFho+YDQzl5g15o3tmX2Jr3dfUZIpTF+LxPQvrMt/gM8dy9b8a3oETxdeOeY
RjFWZFXgO3VPIvjghgbE9bv1d6d9MJrowF1xQBSoH7wHJGJqNB0vOp4BGcH3oY8j
gxr0oAjXuFnkseY/8BAzJgJ/txXJ5sYCa2a2yAN7qME1Rpw7NHEhAzepmdZe1icn
gs039g6gZycgigYq/Vn9e9rbFrlckvxf4am23us2Pdia16mkNZSMZzNnz5bmORHY
K+uR1PUwXYRrWszz9+blyWoatC7AohFLqpPgzw1xRn0zmMOvjY6TQ8yVYmKW9TO8
Ysj215gkteyjQX0biMuqzo4ki97Z/CGIwJ4sZTYiRsh/Hxmo5BjIv081m/eL2coI
OPWdCmnRUOIFqqmohgcmpqrZHzDtV16yFRm8Yx/o+MjZrUHsFrnIifLddFb8QXTz
WwtAsyG6jho92aPL09i9y2nNkSI3db4tGaCS9VHeP9miEFV9S4NgL8B6X6GXNhqy
AyDnhlSyOFPLMrzu5XsH5LwqXnBSE2gXFzo7uwX89Lv/gVpOJsW91z8lLr17H4CK
GZexOsYuGTJkjkQSBMwBycYfMXXOGFEDhZ32goMZ1sDsttqSnGig5+LGfkXSXSFw
w6pLeGf5Tqm89521HjdmSH7xzBqGdF5zkd6QuZ0JDUzV4Z9i9lTkAdwnsUpVXZWX
WFX1z5mmuj2LwsNM4Gtls8JqcvwR+cC6k/p5Yf8hJroPAAKMzO4pr2YgZsVBlnk3
vuauri73VcEnleyBfL1uSCno7F8jQTPqwgnbuaekV2i9XSEw+s2shQ/rXQATZ3Dz
JOZOITtgl2t0SpgKCUyuMuyU9BnmsVcTyOmY3JIh092xV/2KZRLFWr7Htd2u2nwr
MbqPbXCZLF8KRugS0cbU9+hiL3F7JA2RIxByMg8jyYmmv3ZmGwM52TtIaSQtkfok
Y1bryVLr7EUZBncFIG36mxrEcnqZmbpZaC7lxYUFPly25ZWIAV1tcOpoNAxWmvt1
V5TnhZXgRv/2umpm/0czJjp1pBQigtbMrzLQoMih7UCMedGqVjaOuet1CpzWOCwm
QJLs58tpNMm9byV/JjlS9FEmSZXVA9g3fbi656FZ7CODi0OKWe26CaOIES7l142w
VvNdWiTXzT1DdOze0m7lsJk+aVL14xIFwLFy/Dl3wFFDUZbGuSZscg8f0dtXGJXo
a0drSwoKCwKln+QDZEpgJ2wH9OXmdqKbcykTdoGcaXLVGkkuK7EAUnGWyBN5qoUR
rcb3B35xprkliap7nNHvlfojFvWwT3Ki35KV+1gzb4OxS7Csurs2Q0aLIJw3s4E/
LMkZIWtnumNQAs59pt2fxX/e+/PKe3qt1oW66vKt1CywoXUyabGgyhg69XbpJbEM
5dNdNlvFUWgxdYC3TlSGoHrcvPZYM1RaLlZRSD+kclcePqRFCCyWpn1xW7oMfwfE
0LH/t0sBeJqr0FVR9Pv1Ism5MYGmUE+dSyD63UzfR0/IVSYdG2A8JJGozquOtrpu
J1jee6DsYMwXg/2CFZEtlgJc2pRUoHyOn+yyh9hlmOztc1egsY8tUsDQanEXYkhX
JrOFOiQoX41foP1tBw9w1E4hEKNanG/Q5qvsEaUtzwR8Vm99vYFHITs9cMwRIlOe
rrjWiaKli7G05vtXjGHl3GXZB66bAmiXk1O+1PD6qlagdlZVjh7Um17rVvCpq843
AxKBVmXHhqreXfvCAchT5ocpllu/QMdALcGxaTk0tKshDuQgn39nKUhz9DNmjKDZ
69dFcVdutKlIyhhHvE9ju8Qp1qIhJQwCDV/3yVQgCPxmJY0kk9mrU08XkHi4GC4M
MThMZ0OfBIbyb8ubniCwr7jB+fYMoLp+akKHFpnmTHmCa8I+RuDR+/U8dwCmS98b
urkR/MYXvelg4HeZ2jX/Itu6maVd1wSWf13ghUQGwCgpz8t4zNcU+1ZHnKm3bPj0
Meit83kEUI4aQo43K3b4a7WSu+k0HCynk++TK4tRI/8S7St2VZ2MvrLlcKsop0rZ
yReSVMYTvkN5YYViau/AhAW20enXIISQZFQIolzeW/lMk/vBG//Qfibm8hvogkQF
264yry8OZb7ECgI64u4a1O/+TUpI1hOHGt1uUtQ45CCD7DgHVRYeFhUUlo8qEePP
dnPVwrUMQcpHgvxmmjf8DEm8jMAplyAuXv2XpeOqfBTtY54VAZ068iSrYnxMjLAz
JngGJ+ozPpVDGCLFH4UwHFlLswpBzwosAVP9Ta+As+55eRMffdwuuVKxpg+2TCK2
NCiLgPbhAQn7NqRJYuGlkUSxGxQFVwBqwYlWGd+CLdWCZVQX8xiOxRJXyWCuyqZB
RIINBSRfQatOA5ZwJlsjvXut1SbJgJzfu138AG6l0ecWMjXFTbG05/N8ESw66EXf
WODg2zxdsz5BiNNDScWhzpFAAfZ/sosF/vnJKPqWjCavrBDrwj1HMZu4+BIRNii0
sfLZqaLr61ph2PghjuL3QoGbz1bMKAoOTMMXWQiVlRadQSlY8QjoKJvOFqEGkMZq
MbR9p/l02s62uiQ1Xnsmg4paFZF11n0D9abeF5ThFLIFW6jCBsHcCYY9ungMKlyG
fSsLRAT1SIOFtuzdof/+ds/qYPdoGBF2LdqF95zEbDyHD8KnkMvr9LzQSeoF2s9V
aacDRxkoD1oVC67EOQeUsd9KOItugE5+9NhKbAmXI3bR7O/rWOfbBrlP2ADvXwL/
hXZ/F067XGhOSIMLCxaiw+OMeJU3253haK1DrFPqznMe4C8HSxLa+XWi2iJavr0d
rS/K61geU/8KXEBskDun4cyo9REMJpGY3hqKLoDDv9Eni73Bm4mbxYwE5kkZ2vcp
WRz6TI4Y+Zt9K+qoZebfv+hejYhahzt2+Jafh8oAGOS+tHCWkzO4nwCEjvVM9TS2
A2eANw353rRqCrCRzDdXgkFvQn4J6tXqKttsf4acG2wGB1nJA2u05TzEANTn0JWf
7vs3WbCBNzZ8uMxQ+sjQKC+F88zOckL49Ofwkc8Lc5TQqmwFA0KjpD3VyUfCD/H0
UufO+fuMKZivnbkSCTqyJ+VO2ZMlWBBZSfYaqDDcOvemkp5t0uMZtwPV0dDHYurd
U9uNwVUfbJZnh0ojXmLLxOxj3C0SZiJmIYCpNg6artDQBz+S+aXlBK2b2Rq+cZAw
FkcIN9v3gqUxdE4Q9Q+xjePzXneq55VeMwod1F2rSWaP6F36n2mk5P3tTWQT7hnz
khxMzWkJcmtk7jG4kviiFdR6kb6ZU7MqdW/5DxU8DVuOXPA0LwTlmlH1sTEum6zz
1Pq1xNio3+YZodPUL9Lm3ii9i3ISLSRAjAYLdJ9iwS1C0u/mFUqVI9EEOykmwisp
2Hh3DhOiCet7nRe881VtwxRDcjryu5wXY0u8VyCX39Ts94XIElJz/gYdrufghvgJ
OGCWihkbh4nC7Th/jPydl0kSNKga9CXHkJHJchQqzhoe82Y3I6aFcQzuEyAJ1YzD
aR94Wy7VkdVp7IK5wk065FOaLkdU9YVgaDTP1A2qn7nFTalE9xLUOLbufP10Bxi1
A/JLyHhi/Idp08oshwVfn2An/5og70AzmVOvtRt5WEUkEwAIwzTBN6CXbonOebMx
wkWYoQ7Dj8FihYiJPXMDB30h5IBQ3kW/q6nOH1nunXLvY0IOKKXyMXxAxzCaT6xl
4NwTDdH23faF6ovaTgc/iVWmba2t+NK8CQTpwDqIhNmWUvQmDElH99H+ReuFzXUu
wLGJHqxeYwU0wuyDO800ETtIl2fvBPTxTJDEVi2sKODYr1re9kwLXCge5OpU46Xp
YlRpTkHrcvo6UJ2VY0zxN+JGgq395gyTT3kRgzTM/0fcZArc+NYsXRB3nXRu1u7d
vH/F4F5srRL1o11gKXA3BIoVVjwF+Ft50a7SdttVuTli+IR0FHe3d6mWjTQ7KOrH
FDFgKtCnjIoDHBlz1uS9KYlrS8GB1oBd4IRn2grCjaL0IQsfjP+MM9r2irMnBiIw
IBnqllQzW9OMGxKZteyeeCV9C9UxkG8iFpcJz9b3a26RwcSkkQgFRpJxqM27OPmx
PBK/ZDq5LRcV4q70g8DDxpzk2nJ5hGObgvDyvEY4v+z5/lJ+QfkV0laXlQst4Wkc
pYp43yX6IfrIDtHvNwUHOD9WIpelatMQq0K5TLM/yK9ArpWOHo7Qx1TEinNPj7c3
fh8WG7gvbPDrxC78ktR73OXt/R8khe8LI+JN/swvU7uJMJY/nddHhapVXGcci839
+728sI/oSIm9F5hh+MOexQLY7cWf5I0xLriLSFxuIqnYjjGNGxXfxfkVqeuCRwSE
eXJKC+p4ouoWIxV5yMaLvj+3EIoN6qBkWj8O88JQE8gYiWTT6ppGi9AL0OIfmy2Z
GsTBdLuw5sC+R75E7aNE9mCo2e9q3cD/SmBuoT1Ud87P/i0VzN72fmCN/ZjCjwXb
aoEDC53XhET/WKkgO2fQozrBE6Q7j9zSXoIeaxGxsMIx7XHSlbJhkXla+U6XaW7i
smsBDQAqZUTAlSJfKlGVs5OJp8dOWfRmz/+7HA3y40TdY7l0mfOvn1QkjxnA+FXO
svzfXVunDSsrlyZ2FRhum2JVHp0z8vgvcy2eq+jR3zTTT4S1l6bb19EPuPYoG+QW
1MxLxpErv3goDox5d6HPLdGw3numCePfvmoaKncNYU2MOSWQVER5Rc52oPJJ9VYP
qo214/H6n7MVLZkrGhT175kTdEiUSGR/dkQKL7g9JCnVjiROaxUQCMEK12n8oWJ/
nqlT1o0oHJh4fn/4SWeSavPhsjQgXZ3XZm/YDiN37sQk7EuLEFRyUGdsoLQ5GUgL
By7YNPB7WKaxN4ndoPHWB0Tko2pJpA7OjRrBRL9u+0zF0m34leYxtF894RNRsmap
Wqx+zylAnVbUn84z5kV68OSp/v/UpSMV8n8b3ReZR6RjjJComWuhXvBkn9iNdHTi
E5DYPuWZan1oEYqfffzqeGWJjyyigfB98TZUzflSy7nPKR7cOBL/XIJT9HQqmAu+
46+z/CdSHWhKkW6OOYDJapKbhTlEA3GLQIcUHrXYRT0IZ+GY2c2HWkqLPG29hG/L
9fN2x9+CjfDLCigmZcFVZC3aEydjtq0EI1khrkloQ3lMlAuKpIJ1e2o59bnCV9Tl
+xGXSfsiaCnaT3qmFjL/bw+V9bKkd7PxsE488PgzhwvvC3bgUXJdabOMFBb4sTyu
dbc6t8VopzjewSb8+gSJ+2H0gnwtOvJnPkdRKUB5BLlELU+XjXkJkGkPKvfPs+Dm
rRZARlVMqwk8xBCAxZX9Z+4bv9pu/iP3s1Uasy7AJCUg3bS2Pr4K+AoNpSTFMgnh
Z3IpqVnvlBygHqya9JycswvsWlPP+iw+BRVkeTqAYqblWErw81vHmgNh+JDLgB+1
YxZTOR2MmvU5QpKNiKsHzXYL4ZEgBEWto7vL0BHshN1yxjLyfMi+gtWxgOKNjmQ3
f6Q+XeE1ULptR8S6Z5JMxsWPW01x24RQAk1Ji7JsK+eIiCgtJN/+JxHkqeAESWvD
2XEothNIxs3XFBA+6xvX9+X0yUhobhilRO1hmNuU4UdKDcSx4ieMtj2tRxt1ErtY
IjK23GJMcHqcNSQniAZIL5D0ic/WGxXXex2Qu8xDgizn/1L6J9GS+nDfbgZsgk+C
9wPfhGHwwVLqnfhpg9YTbUyVPOPEkLKuhsJBnK4Di/SsMSFG55RWDRPyBxeNyekH
Ond998QUNJJII6pC041BngjKD47sON8ZX8A7jLJa2l/YGvV2Qc/aP8gvnMBykceM
wY/+tdOTN9/d2Lax3/EwWkvYi0PveVBS+JQXgxE6tfh+U1EQQHzK9ChHFuhhc5vo
cb7zLLwTSQwf2DudywyVt3AL7MP8I42qWc4tHjeIXkDRiQdHY8oaJOKLPTsweiuC
/kiAdsqeDWbIt+YO3EZ2/6SCGkZS/O7SXWAE6OplL34njtMlBQGmQoK2GC22+HN6
eCX5w8LnMfZdGWQPylFZHiG9Ho9FFa05kXtgXQ8W+q26nkaffrE4cnAWMJFTKqvo
Byqvl0DN/Z4cZmF0u19tncEmmUP8kV9r8FM+bQ7UGAGcq3H0J9eu1mN3KjEKdDxX
zc0MF6oBAJoFRGVq9KfQwQoXc1fRlQ8LVWM28t0SvVPWpB7GxhL9PSfwqgU2lXfO
daCM0iYhLsBegQGnbuQR+wKIUqdiZ3+IGXCQT65GSpEaoTLI3gcSDbxY3utAGTRm
OZQrJrMXiLPp7CUxyg5GbqTOO5rvjUayx58j+PRAqahIO+RbhuX62VrGbEobrMKP
l6QTwp828wl77yOpUHtV2ppvGLFbzsaR9EUFTwXpxS8fxQFAPpponkrUlZJKiNP9
/I1FuHsGQZeh+o/S27HgWGvStXtYnHV5Tjf1TJwYUB/VHyKtJGCKqJn628CToB77
Zfk3eyH8h0wvUniB3942lBstZAe9uk87Nq71MUpdYMRRoZm8vz+BKdIzpv95W3da
nanbSRDaVHndQEDr2OGPF4e5fCarVPcd8j9qe5bcjGkdZOjKBjGFJc1NPFSOF1AA
W7KXd/xUTT2Vygd5NsRvCn4vWEq6kDVYz1VbNQgbfZwoK7shIFiO3oa55+0EA9OC
QZO3TDL98wfPlPRfcRGCxnw5jQMYvHXGKySoamdc2JNiyIFGFre51IrpxI8x9lGC
bTRi9JGGvtF1Hqfr6JyPf3KCOpNA1nubzprrdaPfkG0NZRTKFM1Ss9vTDZA6bJON
ScmeHUtTqR/H5pzORI7uD8WZd8stMcK7r8aUFTTArhU/cu4YTZE5Z+aJahRixE98
4ca4Qk8EHkLVAk1xSpv2D52OwGc2khGa9gzZNbRy8C3Le4tM3C1X5bEUt7UL6BCF
1w9YjKl3kVmbiSJoqS2Yy3dX1Og3PMZkVd3e+vPtpKjuNHsrm0/LGAGJW7iPN541
TP/4s3lqaYyJ4a55wTiepXLtI+T2K1yNfmnBk+R4UcTJb+zMlWqb2NlPa+cQ9O3o
4aGpEit0xKhG9BliFsYhFw9Hrj/QzlzlmIdW2xW331qYknj5v/WOADc75Ikg1+6y
nVDB5HIhwvdhm3uxoqmSp1lEJNLVU29lQzVyXjyhaFL2EvH/3iCac0STCw2Slcq7
hluNsj6pjIY/K30WE+dC7p7vOtmdSrIAPsS9OdyNLpZoaEIkSZH5bXahnaFecqOk
G6MQo6Dg7e5Hly+oe03sauQvQqsDeglVD6+eRxQcnNXldnpuAd6BysgWTTGXd2QD
4GsLwNQNP3UjQwOfPO4juwRJSV8QhcC/a69JjZbPsvD/e5w1J0njhrUFYIzn6q/p
2BoPBXRJn35r573nQG1QfK2629AIT9lmzz3VA0nSHrY1HGjJVz1oSfheMAW5bvdU
u9HOc9LagPDPMW0oNza0V5th8j6G5yDV7DtNHbOrzRXgnor5Lyc0DnQV3c+RGTfs
bPb1+IQCBTKMeI7C9Kd+idZgI0NUSb5SvBEgoVtdRtr7Qw0MBcEzE/IVj7YHdpPF
7glzQ17Jo9+sPm+rl2Qj8GQLGI4JzHiWYRK6fEX/U/eZVMedCiadssK2PruN4XHg
ShsRYYTdjbc5aGETncQmwRC2W0+o5EZtoFejrPCm8Z5HBCkYlLo2T8Fwu6tP/j+o
FOkY0YRSp1hW3kMrSEmIxWtTOk1ag4fRgLt4Q19DEL5RXG+DDynKFfcfPqJ7KiuY
LDeHTAwDpkMwb1PNYNipSqihKIY7eXgoRTWSNoRdW0q1lXJIxzxI0Pbesm+EYjPA
jgneC6OS1g/s41HGflTZJd/bI7DjsqwBQidNtkCf52EVGaFcFi9eJxry2FLWeUKT
I4QsSAjVyK8gcppF/8NtZb5z2E2d5by2Z29OnMWGRxbZvb6MAvkbPICn2nu7ay/N
xkLBLvEHLit+lPUNm6SuLV7MNQ5A7o6Mh0A/aNtyF+DXYM6RZbqF5KdCzQN8E6tM
au/YYsZPtz2jUoh9OPv85oSCKpHTbAgT5qg+2qJs+gSDhp4ZwankHyDvnLEcSz2n
cXHKJ/fmmPuOLtHaJV+vHAJtodbvELxUs9R3p2sEqujzp70lnY1BiF7XXNF5bfjE
TKe8UVd31+roabf9h7neUjMleFqWY3sZLHnlJfIqdBX6OUGVyY44bwa+iRuV/6Dl
ZX4AbQcZdF8uRd7lAzDrbaBnRC3qyIjot1harCed/UPJ7ryNa/Rnhybn0BtubtSJ
CFwM8tAu6QiMWhtNrnuC8AD9zxFm87vVbQS7duaxxAQ41VtXjbvWXFLykDaQBeXr
KOV33o18Du4/11A/HVGA2UWOX5p2igUUNRGdgGFdi+40Hz6rmqKZABfAsu6Orbly
QTrngHL+CLm1Ah7vmStEfqbcARJNwoAndWIkwL21RaHEuxw680f1HcVzoR161fWi
32XeMp04Bf92ZYKjs7FaKzoYd/vWPQTV7uNVDJEhmoKesmmTKogNkpsqHQrOTiIK
NLtphRFqJLyO4Ay/j+I5dbHE+GJe5wrR26g3QWWkus+c60yGpHh1dPSH59Iby2/8
x2/HJzUtdH79k8zOfMz1fJC2a2sVKgcJqzRrzjV1jZdfplqIcabAqAN+8h8qqfKU
jXEdrbMxBZg8SKGfveO359oPT34tPHlt+NCxDorbdPDuWwVAAOj2U29IA6vbNqBt
vAykWcfJn2AfK+IlGusnNletaoF+MeZJPUR2ryMxUPvgOZA6E78N6j8BTDCIE7kz
nABXrkuomvaa8Uob1WNtSUta1h364a8jFAGD31XgXtJvrC/eMVlerF58cCXXqqH0
y5BvZBFD2niuwth/SK8ITsq5/v+fr53PDtDqecbyMXlSSZ1WPsSy44Gl9jb5085Q
RNwngKAYypapfmoOKFwLRtKiuonAixxAqwUf44k723tAFyQee5trE0l9i68IsnkL
oGGrh/VzWJeLh4ALlxSiV0BzOynE/Zi0NgGeCMY4ItZEGLgIB1C2slTzdC1/jkek
EyavoNNamrcLXhb2PO8xTvXcmkEkVqAU8uf5E2ZKfyyt/xIfjoe0l85H5GOfSgX3
Bwq0K+1HTlwNkE0meiSvoVWsmTOjTt4PMQ0xlaBxgcwYx4PMyVdGZ8oHkWvOzGPt
vapnXdxJMmiVN8UYy1zuOw08tiRy+djFqVD8+8b+KFvpJUzEL0RxvTj9Xz5u2uPT
AJwwODbKcCReYbFPt0TztIZ8NP16/znsccX4xfl4AZEoVzN75RMee1v4J/EZQ0kV
qiRw7TR7WJ0JJAjbzPyHLa6ukUHjhSD2XfR96XhX2HtXTmdMT+ddTRj+UHcV3fg6
l72WBpQHnPDhaDcsxFwADrp7AiGi2uV8BJN/n6KkD1EkcbpMinW+vg4ZH7IizYxm
frxW6L/efDCLzTQbVRxf3uxLr9J7GFZ875AhKr6Zs7mx8GGTPtG4ELKgpFeby0Ja
2gj9l44vfDuoh5+ujY0uxpaSVWmtS3R2mJ4wGrFDGwRGz5BIhijyQ6t6LbKpM9s7
P8hPBzEyd6PDjKwVHQ7VYINYiux1nD1s6uhSultwzgV7ArEtyRWflkjVLRrm0Aac
L/qVDnSs0yqfMzNqduYrc3SRflqh3Q39Dgjw5Z5liiPnWHtkqHZZNn51esI1j5hs
REzOVIzySL/jIamxuBvxhlehAbfvgb7eU1VDiDelxNfQa1Jpl6AZThxbmivBeb8w
jw+iKgM2Ueu/jKrrF6LZ3YhYPEsbPLYWqeTkxIyk6LBMhZLpiH/p7FQAr9id+StY
OxnZMoQRbB1UehuMCEpahKMLgW1O4dRUKfx74xjBbImiWhxjPihNx42GZV6NIKHa
dGUf77cMVCAeVxQjFBWiAWD0lggiGbr4rXp1sT+TJeeINN/3UCMUOmL4YbDLNFa4
XU+ZAwCDAzIhnaVJ0ttMUPjzNzUcuB/s0F4JNonJETFqN9B25QnDXlSIX2YRR3FC
TZeToeSj8SmlAhUDnle5oc3Der6P7KKW2qGN8Id16aHfudqG6RH3HU4G3GY4Jzi/
sHlD5pz0YY2pqcoq9UO84WWnWY4gQ0i+Nph0jT4xDFjv6oebunVN0ZLSH4yyATRv
Cg+hiCoXcCDrYibgX+pSHjHE/4w2ztzczlq8cOmjnb14z7zM2kSZY9pg9vIvXjwr
QuJMnzkzWHRKefV+69eTJ6nM0PXwCGQtWXFYAm3I3r0TyNcdmTGOdJT77S6/XcH+
U/PJgwlwy48rHOZkxuTNZu7JUZyvupnnrVIbz4l1mlIj4psJBLMNtyGjiBYumsbx
tlTqViL7BoKzc3UDrhqJ5tavT2bGkCgvzi9f6WknRBxhr41h5UWd5BwdR2Wa0vw1
KmLzuDOUqn32/D4Vu3veLnGHNcazl0KhGod10d1esgS9+kWSSWwZGuQdckGrosAM
KBJ6uNbbmT++tvPBC4xY5NNA+N0iZfE8wztYlAR+Y29xHMRVmXj5n/29w+r1IxJl
OTzX51L5a55X3v9en5zsFzsmpIW78rd0K5ZRuQ5RK2zUOvEMrxjvT4zMw7aIc6ME
QujgI6hwFq7iocQs3sbHt7HpNglW3mWsgAnHYaFFFQJf1H6sgIN8RcD7Q++R93UJ
NvMys2Q1JhDTM054V91a9k+r37NazfGm5Tsfg/Ibf54P6Sq65fokZr+howeopNvK
frUhseLlaeprVQzmx21hq5zsnSrXUNgAWGG6t/z+LtMf88+bes0kzn7XlcjVdSF4
4Rf30hxEBMR2E7cGK4FEzEu2Sh9MHwSlx0GJ3FbZ5xMnUMFtp238V5foT5ZELJCj
UBZS229+COalFxrg3du7AtAw16tv8wheEdmQ02NZOXNvQncZ6hveBWG+p8+u6G5t
1iDVXVPbbXJe7Z6uNxD8qrGkjs5RoK0Yg/016UR/cXhPnb+/fMyasjj8OB2oBcb1
eFcX1gIWvpbr7yq7u6MCgrZnm8JvKWHnonTDhmYDj1BHCacRol4fuvcHXOi6jHPz
mjU2/Wi1WnDx+qgMmkg4QsHR2PteAzxE8sWcumpKw5OQozI9IoAQMJDB9nGT8c4W
v3ZPPUf0QxcZQqAZOtwZV434Q0tT2Z0ApWCi18F0Uhq1GHB9snfjnE/8/LXSawFr
9Rn/OnjYxNUAsLmVPlNiKiK9Lo1wZ2ard6Rh127GsKECfUG/7/LIk7am2f6goK8o
oI3u+suoYiYq8Uf+QFW1LwddWrjchxYMkPw/30wN5aKzKrTon1KwxKd1HYJSQVKG
zUeO455II+CQpTi4TKgNvz2TMwxffoVuCJN+JMQQFrgrdG3ern3kWxVko2EHa6VL
SkgSh64Pl7wcQCL8p38kXEub41aCD1KAeH7fmVQWqTl9tBtjIxFqZAsM+iZ9//Dc
I2uafjDM3Tr3iF6vX996RqQ568QIkBDdP6/D5aYm3gOubtNgzFX3HGcOA5Hu1yIm
+5xDSHC4VXxzIrxnP76upfCi5qIbEogEpAUxmVqn1JTAzoXXHnfunhaM3KJiZs9I
ztCMe3UWXwJAJX7fkZ9a82gnRY+FYq2OIiOiKg4VRex6CAPT9GHCeZTOhDN79kSS
OduJXxWufl0cBk1VYcDXRG0VqcRNSr3hDlJlvUrW0dKHtY/vOql+KqLZcP0rcO1e
ILHLLbCfCDeF6+5wXT5Ft7pvsztQnD3jHfwlAB9qfgaGLsjSe2maOzKFCZNvNhI9
jtEnd75YcJlbJu5mpTG/PWref5ZAL51twsU1mrMBY17grV17sHpURzGb0WKokx4J
SuY6a5wJa0ntrYONhbhVWZyPro+KTUEshsqoRyy/mfdZl7x4MyoydeXPUr5Qeknu
bukHDsVpUrycEKNRXRJCYrKrBSLfZhV67KkJeS6WudPrpbUEw3d2QPVLQs2pK5HP
0ZsKmBUrLyyYjfbWx5RQcu6WYvIbsvtBOfLJXFcAxlPcWBWUHNkSjJKpAqMjVGEp
sN4wnhr3GIJCZLE6p35JIZkP/VobPkYxkuCAdQuShf0DviJBTnLKpBNCWvFGl5xY
hCc7j+vALdon0PbUxI7O95O59hoFJx5oitc80HhwyceVYVYAC7+2tLG2EihQ8xQy
VRg7lmfkBILHDJH49ekL8koFVA8I9XBcunBuQVCspv9LXDXb+1g8z+awH/e9O54u
rkXiJoXNzGmBlKGPTwYdfeI0b6xu8hCJ8ig4DjvL5KQLn0VLMcBCVo78Xtjcobc9
Gzs6tsprYEakGXsQ82bh0xz0hLEx0FaZJbLAchU8YltvXrnrF6y776I814d2AaHb
yIswIcIL/iClhah5kWM6gAdML+nKupw2oY5SjNdTw0Q3+V8h8/65NDWmmEOOTtav
g5VTqA2Jezpdnr7nLoB7ClkOYShtWb/j/7Qe4P3Hur+58WbNQWMgQWb/6uZPfb6b
PY8l68UEVI/4ExwFLR6I7mmmph3RxlmdluO3wJ/TF9pkIAKx/yffrx2bObHw4BhL
kwZDMrokAy8peUIeW86tSlkOrRvPSdSywRzNzg+ZlKrSyBPQIvGiGZOV4f5Yl4uo
wNz2sBLWcxkNJEkwHbSJmBt0mwfpq3krrNdrxmA+4/8dlIrhXHoarfMFJHya2tTc
GVCa3f9N0wdF4N2Ma9DD7r+jQYot/4ojhboDBIfzmD9IM3Z0kEYaDwCB5L0NUkVf
tIdLm2t+x0IlwPd1eUTSzdD2LfYtXgCCM7OQS2HOGYVBcKXC/sisFmuGQq1DEeRp
SBu12fo8HrUoEPp1BuFrwC5cqiaUJ6YlKFjwe75wIsjUG5lKaxEbscJKmw1uJVjO
IEyEKW+Btf97luwfLh/UaF1STox0LtnebnodHo8IqhKU8Ip2z0ubwLiTnB4eGvqI
aGFXLb0ArgymOHOwb1HCLtQj5KqfZQq4ewxIN1y2bs4sp02jv3PREwFJ8z6YGON0
ofeHIVxFexxeeyRurLQxSF49k5OaN3RQPnw7XIDWDw+LlOi6HYabitN0DpJTlnZ6
oXfO7sz2pHEf/XwQBxxOcf8zNyZE6Jc6o+2a7RO0NkrjTAJZergyL9em8ZZhzJ/u
k+TJ2qat2EakydzQVCOfQw7574icKOpsMN+MqjkVd2lOt1VYqQt1GBFzDYGuhWaj
M5wNDtQ9kPHGGgrQK0o/RL6GDUudT8e4xJMe4/Ybpi+IkandjOHTeBA29N4Y9D93
ki2EkDy154wlndos2kvQiaXA7+mvccTxpBMxcg51GGV1scUqVVmwoWSQY79oIQe3
k8s620CiZmImp7hPEL7t5SHZaMEx3WFccePycJyC8iVP4hJ4chwXk5Q5pFeHkwyr
ORzTXYgwMeRJK4/JZrgdLRqDYgTkV9Zn/8wBGGQO7nzZglsI28LTfFsneX5CTtj6
zaN+QKi3WJJOjuU/vFXdjb1/DgflqJqe4hYQmzgrGrCbcW9S8MAqjOGLZodeIifZ
/8d5Mr3XD2tV1VkHuq/yOx5sR1+FVV3riXJPEh97j//YimiKkTLFldFSd+H9SYUN
C7Ao5emhaigS6tZbuphhgmAgpCZBemyHE4ZCWIMn5OEBTeE2fHTH4x5Hv2NlGJyy
mvbY6z3Fbfd61RiuFBVN5fqjB2nqBFX7z1sbRx+MZO9fcbAOmYqmyg37gK4K1MoG
AH4VBG/4obckoNmJqb90Z9OEU/oUOQ5+JWc8HGfnNThx1mylPu4wtx+1P43kYCZu
pRXql7bFn0twvEd4B8YFH4WbMUz3dwUp4yGex1FRqBLPYowObW55kMAZgo8dw3ih
94vMAJ7LmKRi2Uc2b3gKMFXT2XM9WPkbMytq0NN1uqegBtl8nbYljP8bejuXkvlZ
Bv+PhGQyWrsecttlSSfUE5MlGeYheWytxl69BWfJa5T9/upWSun+jduxRQKZ1lei
KfRhNXvQKqQJ4CqXOpIZdLt24EuCT7DRhvnF2olu4YgXAv7bS3kfVA8DjOCdlYxJ
Au2jzLbeIWlnDDtsipbceoNrUeu/DwgeGHjTtypYoeftjdZkVzPuKgwYUMkz6YwS
jFQRwrBBw9gSsl+PfGzmXRzQn4K/PWZiCfBpB/fwQ9frjAq6ea5l5G9S2OKam0sx
VXjh0250xqPOzDPhW83YK2+Tk6kMh46RU8ITooauve6JkivgnExg32KEhIQNHcpM
95KKGLf4UCxfYVcxR+q3p3eT/nq7Q8zBZg08x6T9dv2ROnGSIUR6hLaLQAFqpHAs
sjsSPZJ8Eh+INkIuHgE8etoNuwyKROri7E9eZGOBNpQW5h7wVgiM85pUc2/OungA
ma8xiFjbPMlbUOs0FAejF/QVcYBD6CNFVNu+IecuQ+zXL3QugQLlBPIkPHGmX0K7
rVx9HwmKi8lbDXQUZza7j/3ulR7LQnZnie/l60nUD1uB4dCPDe8Te2xDAQ0DiQng
bow0VVyOaJUxDMixgAvKAu8sBX1ij+/yWHWZZKK4VE355IEbrtSjlIqAkkRmqN1B
V+CcxouQn57A+zG3LpyBWaRI0nsC6IbmaBHaCm6NUAqJ4o6/qOf7Vf+cfO8njoZL
zeRuosVMRYQrTtR0/hogbDdOEXphE33/zV5jHxVELXJomOWt7PMqYRrkztECCSiU
Bt83wcdNb01jJ3dc8pYnp1gmfnZfBDvoyhZ/nw4PTqUZfcPsDFMi/LI42u1CjTXO
Vmq5mSlvUT/8/yX8pb6jQQQNihAIUtLWPxhCKcnyMkwMs79gGReOZ16E25k9/dUL
/Y76dB1BeSGKUsf1MVZDUkDXch70FK8VE+g+uW7M1RO16cnWPN+yuUZGakbx9LFs
5u3/y8ZjcBFx3Zur9JVJ6AGPX7aVnDdxjq9fVDipcH5XbgXtOVvtOGAJy/vmsR/W
p6+qY1a4AXgt28/aLtrEJg1XjYJ7hOe6rmKY90FhJe0e7ftLaWExyeADJkgDwQb4
9iNHNI5y+qNCV4I5MvclmCAjKL3wNauqGpVcU1fUloQKYS/BIgQZXUe9/juP6iEk
ffFfUUkzSvIPrprJPaeDzfC2q3TYidBkuWgmwYtv0yJtJya+UqQvzFb7dD8hvqHN
elfuQcmwRtoJAYSYSi4f2+adMc3kRFiORqio08BJxpP4eSmiiDqWpyMPZoaho782
CpzT3raBMCu4S90E8jH6yB+4LB/d91weYdZ+J93QF+ciZgq3YOT6ZZxJ9l2IdzSy
tq6GSL8JOcmg9Esqig8D7RzHI/RWNL4my4o99/l/ZpOekIEogj+GF7FB1tVvNkw1
l56x5b7u43r5bB09rL7WxZyMA8VUVNismFcWdI59TxQuaD82NJPqIbcVDje2a12z
7vmIKBIYUk9TlWYS2NyTUFGWj1lLl5JIYa9kt0s5B2M9c5iExEAjoLrj5wLesT9+
vbvies1x4+LfyRM+l2U4EzHg7NfrUzb1hyqjaJJL9o2iFTDa/VyH3FV3L1MoRYYU
WTJn0Etdw96WUVHhvmzaaysSNYYYKR1cfRxri07KHkHvfAFNlc3C/es/O0L0GwW7
f7LGWSp2LFZqt+o2ZTvygaKV8RJWih3O5PtUYEWQsk5RdOJLnrpAR3dBzKAsVRlZ
Hqb/X5A7zl36cY/0/ovJoa63M9bUWPYXpD9Dkg4zZ/OENhojezgSN6Of507YKx3n
H8rf2zX5sFx458KpkT7R9HYPmDxg7pgZ6ZjwvaRUtBjDSzFFHzzB0mPPYpcHSh7r
igdBx3GGlN0eXVaSmfYfNEiKAnT9lQjfeETM2xdC97uxCy6F+adO5Aj99r9MbQIy
QyUpR7ycvOV1d++d5t34Xs9D8ka8nHuXdU7+6KyertRXfpn5BqX568AIHur61scQ
lMF4F+Z6gJvmqqwQC396bLBtWkidkEJRUraKWE4m/nDUo2cdurhd6r1bZSopZMJT
ZqTxulMocrZcoC5BPE3LANf9palrjRCxj2f/P4ESuk48+73hOhgRw4dI9yP+m5So
bHTjOWK1V3zVQ1j9Y08PJMGuinoiv/5scrEvDOuibduDr12i42U6HnkO37s65yWw
WmsbPEgaAEIxqXdoKYQkoZ06b9xD4mmcBP6hjGL6R6oz7fNwtqfc4fgkQlJebUH+
Ay6U5CcX1bbt2Kd40k7m5sLu0Dcfk1vz28Dcx9r3paQUlIp63qeoQpEUniaSBWjm
DygAwUJZVoUh6k9XdGmxsQYZqx9t77L3dUTKLx6krgQQ5/ca9O/hbGPB0xw6F+q4
3Y8Jj09kklcm/ZjImfO05aDgDmm9amn6n9IHy9pUUMjF3+ag8hf2b3bSxkLpTHvG
6k/LLxT3oM3I4gvToDJ1iVHgxCv3r5WBMxyim5eol8hBKgIenbD6LTpZKHcbbPSx
4d7rnBJn2p+e2epYMM6Zil6z9wQVjMg0jBbuio46fcWx9ki9jENtkbChkHVNZeiR
QarRk/U60iNxKA2QS2H9TWq9+GU6eXFFBn1tx4aWgQ7L0/PJmQsHKRGFJCvuDUI6
d29e/z9zfo0A38pAgAIcniPrvw6Dwm02VcJPB7lSGWtD6Iq0gTnwiUClYUqhH2cd
yZomp7T7O6FMJwytxSYxvnBQ140Si/jrEDaDuN0o5nXziFTb5PbNwSTrYjNfJfQU
EFMCeuv4lMkSw5UIAyII/YjnfSxE1NECqwo86i8C0wsbSrjXeD8JeL3CCHT2Gog0
tcWZZcx3MXgPsut8fSDOFCX1CJhBfpofS6fGTqoMRphhL1rEYVLj6TWJRnYwKKG3
fiEMZn2XR+Hr3YWGQFxwahWnzkpH6i/MkGkyz18ohXltCK+o1Tn5i8Lc0kH1/h4x
vSfugcJCU6xW9MQwlvDRjpgiq3sn29xvialmYOIBSPD29C04B3XnSjlA6hw2qgga
jTdWVMnuu7CSXmfbksw0t91Ra4NWaAFTley2oqm3lmKG+tBGIysMdArXnyWXonlp
ZNZaO1C3sPF0PY8852i+do5wjw2ADPyaTMd1//qlm4y8/uCByXnMfK09uGYMrHwe
Vvx2rCgOd2yB3ZAKY1Kq6I2/Y1nxdc9WPZeFl8Fxw3JKjhAH+GMbIzT6NS3M0HSK
N8v0+mJgYiOJXuP0IMtMjHtE+ZOqw94WrMrJ/vsPAXz6STIzyNcQ5gXlJAXx13pM
lqdTIItzoIM6GAk4lD7k+OTaPPDY4ayOwtL6qefSD6iUYC4ZxlAKeAM3JXoPHbKA
qXqQt8dvcvzpCD96trBjCQ9NbXSFJQsJDULn+6ihdUhFT9j/z+QsJzfMcQ7J1a0S
wXuvEg2Hjsf0yuPA2+rfuAcUMIu9/2+FXixFPi4L5q6FQcUGmP8SolNWoaVQWnNn
op4ajxNSfiDyvF8qBy1u39kVoTBCNSJ9P5L7fsXp69w2eZ9A0TJDQLzyLRWEDZ9g
wmBqQ2lM6QAAaiP8SU1nj7Qc4F6X5H8dx6Mi1YfawJ88tnJfEZ3E8RAcJ70kChXd
XiigBvTqQBEgy9NHBY3ITrhLFYfI5BwTLZE6G/DWbzlZ1S6dNEqx3SAhk3Z6mDG2
SQBy7ugUFkHAeyjTy4JDBQhuHRbKdHY/lw9PedYDAjhS9c3Pv3A8PSJM185xHq+F
WPu5rb1UK0CbirZrtkb4XJJidpwpkOzbq1vxzutEKBo4qkYx2nYj6zjd82AI9IaX
tRyAUWEO37LlonQtomsgdl7QvtgefE5+8ImHgN3e2BwBVR8Ye18set8WO/jTzTbr
gjRzqd0d5OKb5tuZd+nhA63o69bfIMFcAoik1K4JKH5O/5af4RcAsuaX/AYLc9J+
ZcttQEM/6zu13GCzBPtzQcDzkkuhfzEpp2VwnYT8xCqrYSIPiWyISRX4JQfv6Z1m
htLCab0G1gQSy/6CRFd8gaGncO+LzoqBI7M5tstXkp5Xy5BHTsA/1bWOr+vdBfkY
lAXlDKA52SQjow52P32EpYihF6FoWhJ4dWyNMth5EpxFUoFKUT8bRFM/ElU3jjXk
t26GPMtRKoubIkigW3vl6iOKqinXgMMhivbOQON0nAFYBPUTRvzt6ipIEz6s+EQk
2TjE1dpsxc8RMh7XQXlMu2T8QBEbA6VAvHTQf9xNgZy/NoIqS2zXZwAx57DNIudk
jry38vRmInfF6o8iPxRpHSzJ/bXB0+zgl0fq3nHw02i4/KCkNEyUFs0l5aIqbjZF
4mopkxDpmakUyWih2QvywxpcxLJwJnXCb3X9SzstDKuBRFP9YDNY/FqTQNtdUT9r
fukVTelwS01OAl2aeuncuTDmeo/Jf+YwoSwvBNKXI1og69K4jIewcGk/iwschdZv
v70BBLMY49aN2eK5FItspa1ZBw8L28h9kgpXMMDCfJBfag3cZWWY/X+TjFjHj172
2k6+CjQ9+pqanJjQgZzIaqo3fo1Kq12hEr3+YaHdtDqwwqDQHivUM0tJBmQeNE+p
VFGz/+AiYjd3KKcmIMlTvMm/b1C/RaLUwXe+L3GmsKSoylCvWdbpWJRan77wOSz1
HeOQ79WNWw7SZ1oI09U5cYNOuEP6pc1waEii3IFoXwKzGO49LaC3T6YGlvD/sZgJ
fjTfxklMZM9NAIDOX30r4ZXhI8eMGWLHueH1dBOkenx6zCKjqOTpKfwhj6xYvAsv
xszOMAGqQSpQOmjGAcsekZcrgjoxMKsnGv6olorrYJY8sua5eiQ/dgi4rbi6f5A8
rNbTLICEbjbzwmUbwL/8VM11WK9d+9ptyaSVgPMRsXgvI9Q7VgKYdiQPISy01+Xw
X7+R7TmjFK/3eod2VIdwpze7Z9HfCA73pr1YjS6q+HBfio7LvxSUbp3u7ZFcR1WV
oiLFasHN20fcX0CungZa4/WmeY/9PwHvT3iQe862h+XibN3vhCBqCqUCbD1C0Rb0
N7577EY9mlKZeewGaOC3vnQDBkuW2+6q0StIygOOlvG8fLPL2HMwJEFgvdcJts6j
CDclNjCw9azi9UZ7tgDZwmV+p6y17utC2zgZB0Zy3cX2HO1SUJw4z0bk/kksn0kt
0fytrc4K81Amqt8aiq/FOjMw7Sj6XNj/svEDSHykTXBmPNVtBFB4E8ZZljkL98p/
4PKn2Ao+mENguxxVR6KSsxFyDrosONeXmrnFxQf9CUJk29/fgTmWJy/ixI0W+Sm1
/lfn+QCjmtrU6+BhKA30IPk+hNkyof+lWnBhceoGj7e7521vGOSRB7ZeYSLfkqhM
5JUYl/oWpXsj/CC+IYuuQ/8FbVzc52Rlvxqm3GY/mcJkNPL+gugHJmY//5kSh3t5
jH1Zg+skTbq2YH9PEMOylWoTVq86qrh6J6XbxS6LqtZ+edMxw+b4wbo1scnq0FYi
jSRROszb0zpikS1DbSX0An9jHqLaTVR/Trzg/FwOnJEPgTyhnw4NKRjubUD4/g1m
Mr+IOyUraq7L5YiEBexwk1DCl9EC6zzbxZpaMveISEIc1DdkQCWUYJ6gvY9z9TuF
EoMnTSGwq0qv0C7f/uPgp05BntW6edQcv/VQUdml0aWks3Xmu+FaanlARbAtjhLT
FJFBWJPwamUUahTkIdCqKSEWYxWgdVXE41agvz2pNC4S+RMswm4REqAa8xqB9GsT
Kb4BQ0+ME4W0RkkFZiXCO9cHWs4SsMojseLc7HvlFKm4guf88//wDax4Q2UM0SOR
pDqntIdm/XB4F5feUOr2Crga5ubNSnUm4GgcjUVLdHHnNbSKF1aiQR2C0zchOPcy
8jBIFVgtRO6g6Cbye99Em35OTf2Ac4FIH7a2KYJ/pidan01i7bRmpN+LNxl6yOvG
x1H9wycANY8rTHvehXmpFAxolN3RxYsAAA5cz14l06aW6piEgJkvhjYj4u94uu67
UN5GD8v57LrsUFhJtwv0Wc/fOjY3W+1yKWztiVW1Hk9ellK5i+cLcTWsyCVQ/oet
+3PLBgzHK3/rZPWjgpp3RqcTTROZShsTKC76ZWc10Etgigq6aEMfAhMYv2k/seLH
WNVXh4J58Kpe7p7N2lv9L+leyeKWrX59qpBRHW6Ss345aryHOpCKMGYY0ijGRZ0j
6BKxe9N8EkroABBtuh4FUtXnzTxSWQKMO64y+lCXl+kMtq3gKE5uZZrqElWawL+N
GnvXEi8TNfRn+RN/FUI6Do22xuVr1mhc3LB6QU0XDAAFnTt390fPcn2f3JbXVSTi
Fj/aJfLiLP1ivGtXRzWZiiKdA1rJYcGjoaM/dV4TE01HBAaZunCCKxAC8knaWUtJ
xQTGFC58PsasWiXyj2hn3z1Wiw7VmhVUNfrlCvpJtFy//I4EMeFWnQH1A2U2oxfu
IWvOpmwUhNtxlbgFVujbLHI6f/Q2SHTBTBEP5EHuW/kH2nws/2jXAaIweEAmKQzg
hQn84HM98q/4TNJMg0BepzDIharq+Uozv+JkvuZAy6QoljouziA7hyX9em+KybKy
DZdV37jtOiqTVD0gOASl0Pt5jPNw4Ex0m6EJJ7AnhEUEvlScrerYtS59/RM6ycwb
lqSKpT7RwTfcBT/vs47FCH9JNBSe+mYxJpf//D8Aya48bGszDYpJKScUJtAoAGF/
qhKilWIYx2syvwOarTVBFRf1sq4+U02t03wj2CRETykQauYNlNsnMzgZUrss+ce5
E8wHab14L0VvjpSukppjtUjxKTXypo18yCpiyjcSw72la5ZNkNZirR6jCrbyPmCQ
8/K5GG6q7FgPYzj3eTU9zXF70g+OV1GpKhxiaMej+hF/VwmqJszmkAmxxcLwVI84
Np89JrxnudEfHK12wIXNOCfOxDaqGDoKnclhPiG/phHd3CrHEIqbnNT43au03kKj
BhI7d+Zsa3SKUZ+WaCHhBGgGR26N6mXoup4hftNYl9LYlxN0T/un/iKlWnnJmckp
kDXfEo/7gNk07HrTmXqUEZllZMhXRbC+ag6o6loVPueGWc4TFU5cokuVK9uZF5mf
bIlxvRb8aW5Q16UBDgwEiB0V59+HXsPnsJc8VNiHzHHQm7FOx4viNUzPo93JNu+/
FCVdy+ocCmDQzxJCyjpHxvyPQsMY+Gg0tHQl0GI0NBKWtvyrzduoGi/u4C0uYjDc
jHHG0MOFcgu4vS9LQMyZmHi6NldtKXLewj0TeYARXnx+MHlLdPDn6a/FwPG69cMO
dn9gYNBcpXv2SjBmfdPalMbewGqnyP1DSYxxqcEM6DTuSff1Qg/XQHzASQrO29gF
UzMLWfuWN7SJA2ss8lKzlA36rLNlsXZJXHVHWZDO+cgS36c6y6OwW2YZIFPLZW7L
t1ytyi82H8uXY9aAKYbNcHHVgsX8dLi+66aRf1ELjdgoAw0uhNhGXqJOwhtt10uC
3r065mU4UhM35ORUj4i1Ewzwj+s1ISNMMlf05MhabDLb8EhjohiRmkzsuerHktwF
GIIdHNsUKuYVmV4u4MaOPmzNCT38i005SQA+dCyUKWQCPjeo1Cmr2oB5flRvNfwJ
FNlD36R9ejo/qXgBcXPCOgEbgBKRkDZv4sH/n6nZWwzCKjSJUTtt7+InYvJfFSAF
kNcoqX+TcGxxkMsoI8aB+7uaPJTj/G9qgGO4mc+IEQMPYi5H5lPNIR/mSNx6MPwV
Q/HLCFt5D/ELTpy9tzKi/Ku1n1W1xfbAM5PUdpLzdySl/aKg87LO6bxEDuZD5EYx
/AIAXkMv35kLfc/Rp9Pdtv00e1BfcK5kOnbrCf6gMbP2ZTGozlCxgcieR53R5s6h
O/LesWRbcTGSGXuv5ITnfZ4AtTQtdxNVhUoPc0apee/WDcHP2j+GmzoxlePz4J5b
05xR9cgmvrBGjg9e/Xzlp2p8LHn2TYVhYYxyvUW0ORp0sag04ZfNmudoskbHa8aU
3p8sNlRi+40uJ9DJvE4+fEB4H4DB1ozD19OF8gp7HKnLirCxqraxOXxx2s4iH2K7
dR7oN9tZ4ZO2h4fONXspd5AceTKXI6OasVrAL4PKuHpFAuzC5qI5Awdo5UIWlR8F
i56vQMqd9uc/6/DQOuNQXCAfH+wrb22VDjE5g7h8mdJt3ZHnnzrUsoXh64EOYe7E
oE3QxL3/1AgjVWT3aKwq8l341YI3wrcIQwzfFBMpyR60dEpXdBJAIO+96b8+qB4f
OEvs/WbG6Ec1NJPYSOXcIWG9Ejp8vGlyIY+KjwCc2wFJVpFqLcFslQvhVe5AZcz5
WNVGc5kQdHdNoCXrKOO+KU/FxjaYqARVdABkRIKB5aoECb/IGtoloqumyjXcwWsV
Lj2ZpSBqwWqtdIw/OhcGDJlET3D99FUVK/SG9m/88gThGD/V87HupFHevA8C1fO2
s7W7ul4VbW464zSlhgD424xM9vDHo3pS3uwZxzcTUktMVjpzWZK1PDYvLVodiR9z
QD2HggspYpnMLZ6kk9mhOl9nFAH1LPA5qcwTh85HQk5U3rKLQcLfSry5t4d+REWn
qPpEPqpUE0fK/bYgaxRf5GgVs5+x1+3PAW1/cgKgWTu3k4u9LSJwE89yB3AyyzUz
9VQD2ehzQs5P+PyVJ94UX7kzO0nYUC1zCm0Dto7QRn49aVvwWVwbhWxckD7T2xxP
aeeNrPBo9oFkhjBxVYtmiDk8xumUYzObuHRjlijtW04UeLZa3w/D6YM3EdEKm8up
435WL4EBgALwkDbKY/RddmTd/7aG4Cc3uvLpuhBKl3Am5F9H8xhCgxCvUBt/ErKI
9mxiSOv9kAj0lA5f+e9sey6iN2vdXZ2YLja8mrR0FwPgzOgPzweSA6wzIHLDVhh1
lyqaMCd92oIVmSqxMczl6VznoksMvHKn1bgs//L14QVeoQ5h8Y+QYjRjOFRUCep6
/qVn33LUMa6B2Vmp60XntAN9wWjlHr9kWXlhnPWKsAVdbxWgbCzEdGCInvfoygS0
Na7w5kAO+9aQiOGQmhWfFk3xb8OaZjZN/ru+YZ9xBtszxnZmY/BJWEi/7wojKOVk
y/zu3DrXFulwZOzWSosH8LzR8gzUTixwxYM0x4Vjud0KedVLR6hlfU9AefidpE2l
lHmi+F1p0hE5WtYY9A2biotrxY2WqbjlXIZNWdIM7gMaE5kw86awGwrLTt6j3RFB
vnJDNzZpxO3/p6jEfm4zhiXYWFLMQ4RdMPuetkq4SPplEtn5ErYGWSe35IBDmyJz
Ekc3PFLAS+jCJuumJ2w6o7Tlx8v0Czv57KfYfYBmyzAuz8oLiCv+dhZY4yf3dlHe
zRA9W3aPZISk5HzZVcVEXCSHh3RQbpAAQ1FGnf8a0foKzHS8POcZqzWWgd95AwNJ
9TKuqywzMHkexKikpn32YPmM7Dxv95YkQmssmTKw5ygUaqzeZxwZI2/FRtLSEtMy
6WhyYL4A2DFEUmq+kTiDPY1FeMGwdRCZ4CW5W9lM2Q0o8wyp/BBMmNJrWuxzQRwM
zB/kvGOMpZrtcEN9EqkR+OYNJ3knfGQ8V9VsmrA4KDhAYvyf5cjCphe9H/4j3zqi
ABpEsF2KVLBp5C2cSkRUnm4pHNP8fclIVw9SnLODlIet1mA/3LlqOWW5OYrPZrUA
4mjMczyTSn7CGJn26ZtcNnRsVDAWU+ff264JayFadh3WLsO5uECuq6loK60Res/x
3JJB48gLivPsebxJnHECNA5ydpiuHbnxk1/28vS4XwXUlau693hsLdbpazcdNegE
wz/cGWCedY+33f4WnODHcKXmNXOCq31aGRBh/uZoCCcx2V8jHcYb9Xrve0yXScXa
TbUjd3fUsRqqFVYjMLQDQ9mHeoAe6UvJ74DizhsFNRxN6nUzwv3kpRULqmavxcKO
lc/NGT+x+nnBpMw7WDfW4U0tFpl3pZKN6MO84I+ovLovcvRiEw4S9f118dIZtwOn
OO/b4JH0gmgm0a8HL+U63fchnA2sSC3HaSEI4kzSvd4LJ/5cvMRYIgzcGGWW7Y6u
1HfzAsQZG4uYxftMsx2hiJQ5ulwh3PQzLGMW38K5c119cyQhj4LrySvP5MczY+z/
NJRCSMrLJDSeL2DDl9dx5yz/T9U1INhI0+0djhuO2nR/g4wjZuR26ZPYEd/xJDca
SO7nostz32yzj9x94JeuRSO7LKYsZmr5QF0aESEha+OvO4CndQgoIGlPKHOIbUJn
somL5nJ/9y8xtK0S8ydZYoyh0fv+NHmgxqBkFOZJ9vY8kXFQ5DflYLrmJgVGpjFY
1MJGVW8ftbMcrSSKTmyzW8GSRYIiqDN602swrMTLs+CmsVsipTXtLLCZhiYGfYx9
7hzAjx9p5O/AwZVpK5BbHJjjwNlOgV8pOIXOYZ5QRQzOrinsZs51Ff+TcDlpMbiD
omkQfpXuE8kWTsrFwm7xPcr4fBwM0WHH1p+dKfMjK4Zf8WxypNPatWMYafHcjvnG
pEDx5VGZQzQXi8lsVM7Cv8pHF/AmWP+TetkWn7E2tgHvy/7dB+bQn7NbqwkQjQyB
Jsx9hhpa4NGwyGGv06TZG+NKjw/yn5Vp70Cj/sym20Re1IpgyZpN+Vnb1qHbpjuy
gcpg4g3iJ1vSCXHz1odJAOGq2rJ1ic2TyyPC0yfqz9JpKUrAymB8W4TMUy4TGDJw
D0UJEiAQ4RMUyY3N1LMKgoiF9CaqKmGUJohieY3C5ISh+fCTTbejn5lzVBKcOn6K
nzP7P4ylEN9s4eFQhqBkzvCEclsr4LE7l8C5kchuplgWg+fuywM+rTGXiFGDU88Q
h0366umixXp8N/AmMeeorMHiGC1UgVhC/FMp6MQvfl38QDbNgs7L2zrfUUkLKFwc
zBf0kt0QFLaz/uCK60zV83eBOo6PvqqlXYqgYZOUUWQUms9vUUB36ZWFpNX+tNmi
2h5xL9EUPXw44LDfxbVVxVUbHOQbULAFbYOAgPeZNvLBdkbBrO5Z/6eZazKCd5nE
3Pq6deIca1kT8yIOvgjYw8eG/FjyyMqhMh+/37MDO8LWd2vslQ+zfOUJHmUFGFJO
cH8PZVlLRAJIURoCkFhXl53ztAhl5LBg0ezKSiiAqjQ4uKcJDN3oV+ska8OhENWe
bFrUqUpvUdjZ+BenPJQYazThKS/aErv8ZsG7FMCcloYL0VhJ7WwC/hiX4MTop+kx
yhBqEnYTJI5dkX4BEWiG99xmYEyWcSSnmDigB3kQfTOv6MjZkfyWcIsZvbsf8jU0
+bwypmoY1sYQ5G1p1po7NXZSwMuQiHnWUKsX2ygc81NEve103Q5YH2GNR6peexXi
5A1J070dlPHWx0GwL3FEI8FUMq+UiRjU2ssVxKIjn5eClmJOi7xKE1V80UAEsJVr
Cuj7F70Jr5jCN1bhhel50q4qs+kNwnaXGqQZy4lazsZ/N+Cz2twhQBqHvr3U4cF9
A3sRU6zX1MFC2C5KKBnKMu/1+7hdn85d4BFcHan8XUEC8HwcjuRn1cOthTJOTIi9
lKM+Kfrk9Ocuws2WCWRdNqBmgTnAD24bRq7KtDSDTnRC+yY2omP3x2MALOM940WB
P07z3fN2Vrhc73rPKS/ggfDoaEiBO62oExNzHCAIcxVndDJojEQpWVbyu/cMiTGs
Dd/a+JNLt8OqJ6A2HPlwjtLWdL6nSn7bw9PYVtgINrvK2nGqTfzBWEvrln7u4wuA
PjlOFVe796WyqpddmqLYACQz7m9+zasqZ+TqqYEbVQfhzMmN0HlvF/9BLGyMXmMk
6VXP3ilKI9KiL3B3Ii5tH15zu1IRGK1X4Y5liYBZDKv34D7lW2WsVVt87wBGV8eO
g+7O/pliSiLZtF/dwcGD1x9TuJYokvLiHp+wmgi6sB/IHKSbU9grqY9pv1rp3LA/
dBC8vK2je2TLGtAN0wBAH7CbLx0r7WIFSO+pO5wrY2GLPMNnhrnf8dzqL6zZgHGo
3/blBeTTP5DqwS074ccOXWkafO7PHUjdDu9P+USl12x2rxjgvdWQJfF0Kr91pUyQ
ujllznZ3UypgWzRpF01bqOLR7ma862jlgx8+ZP0XS2jjy85iAoRpe76N4OhCBELp
/jcnUrT1TxkTyZeOk2gqjQwBqzqAcRHoat5v1jQhXeyfOTzI54Iw+bSmJBFb8bD9
7rrVzdBjZAQqw25p1zGApum6hrcRKiLs7kQXaKz5RxR0Ya5hazm3GDzqBU53Xa6k
v5FkpqyIV4sE51WHTBocyVrDg/cZNgNuQmCaCvVsoMI6iN434N/dof+U3eEksqVj
jKMW4u7Ak4nRKwT4F54/8zEvYGPncgUHEgHWZreexszoseR1Ut+2WfWoQNVAN2gq
viITO1+rZA/ToF2OS1sITzyoy5aiFyJ/uv96Da1bZ5DClELYsffV4RZiTICRiHft
CuysG6SsTWqDzlwR0WoevsetTiUIT8IXbfQuDT/HEGBfSMFkCzJL0krvq8YaFAZO
aAKKDNJ/whrrJPTEf04Ivmg2bkY1+yZCpXAuVv7foKqe+VjjZtrEGXk89DbODWwu
pPitV3FidHbhwRLG8hVIb+x4PKKT4hNB6ba34o+62s98UdDF9x19NmvVqkumHsVz
pRHdTtTHUrKi4e5ky2WmvZCMs2Qrj/+s//5KiOBXTLididiZZl7KogwdiF1G+El+
g6fGtOeFSeDBiNeJslCKilwRCBMLB8saYRlQ//5navV/5UOWeDBCzV8K7a8YRU3l
6e8ccqWs5YZspLimOogp//vDa2rUsLPiDuDrXIjnfabhfgDGF/P9uaLG2yIozXBS
73R21vHqy4WvRfe58NDWgrL6T81F73dqX8nqxiDr/o9Nrb9LeDa9ptxY0h2EjbxK
6VgJv2pMkjUgQv2ciFxHZnOIYj+QT1U+TMy7Qk8kVNaevO9f8AIxreJHEvRsXHvE
HVA61uEYvLEntDsTcTUtbNh7y1t+JlHZ1LgQ9YwmTFkAQTS9fT4WQ8qSmPzmChhk
7EqakKO5mns0v1zzxdqfX9UIZFb7VrwGvknqYUE4D+6TTpZBP1bimY8Di7f7K5fk
bK4Fdg7C8FIx3DgK8rp2mqVqvXbTwKKlkGvYADJbjSjIHSqXPe7ziQxKJL9HdbJn
NN6f1/4Uw4UI5w3PfdxJ8iZWIlhstoCCZFE/3s3MswcYeOJhgy2s5dgexIKh875w
51f7LG7eRxsHvKpJ/EvgvGbveuMCocztMCVvbNKi+XTq7eGqwJT1wSoNuVMpl41v
OADI6BdETDxwbj3WkgTEslhcJHwOqYQuAgdEs88O+hrK10vNLUGAnf+PW+cuXnKZ
5QnfMy6bFo3R9w5v8Bg1qptbpqvX15VtJ68uhtYU7k2XniJrX0JmRLoSVLDDKiCJ
x9UmWv/QPoY8+1YAIuSANhgrCWVh0reqHHa6V5GEzsJ9dDB73bIju5mkabYK1SoG
FquVoRYQQAwXLXUGNcEp4JtGiK7lQxLfr25x7D+VfZ6Qo3vktmlgscOHRrePdzwP
ctHXlUyDcFpt2bj80aPZsWX7AAqzbgutuu4vIFWkBSMZvJJUAmcsFwtXkRuJRgOT
6EaZnfDEhlpZP7eUadMEa2dchhoorf73EEH/a5JbpcbpyOTsGU9KqgGqCJ7KqBJv
31pD8Z+ytcBLfhy1UhrLT5ic1H6/n7qJ13dUqGt33/fRQv/xMFVNw+QoLQbbHnGB
RIPAfrsqHJaeSe+btY86E1pI2CCN3DoTgv1uWjTT6mZQMWkkFt2HDM/s28FHA7yy
kPb/Oqxz8LmvRtEazk7eX8qe8P3LNddGgS6rPsa3uKU4hNucIbcX3WspItWauvzk
Rz7cjyiibUIRLqO5vZLmWrAqZi3qtnysIlBbZcWw6rqCBPnwlmvjKwgfm/3nuR5S
uP8KK3qSImiZsPed1W+hoOTe3hlbJho19jdrTZ7bd+J6ivg3K0yxgYW7vidSTskk
H2XDixg/hFnHRdDn5cSCJz/ELho4+2J5mQ2wIWJXx0QKnDA/LsW7yikr7rzEAqTT
QnOkC5kUy7TL3nlhm+UH8b3HMYNTZQntk4Y01gccXa1XP9zv/B9ogK/08g3xxv9d
BFVhT1k9bwcKlQfyaBhrNert5aupMtocTkTaT/61EZtTRotM9nDbYcA+w5ss76aN
bsw3W8oVoLRkc1yw5p9Qkdl9Dd6ZhUnWj3IfY8xXzwVwcLnKGe11NDcvh1wzav9+
ovc9Er/nHIQhw8fA7TnyE/VMEibaVQFaOIq94XxEuLZWUxQDKYio1xu5seiSYmK0
BvsqH4zT7tYdQ5DxuUrg6c7TDWM6hNT5zopGN4WuWYNQGk5iQuC4WAcZkyXGSSXf
KyEQb2JWYFfZyRbMDqyZPLDWl38u/68mdzQ6wVNmTQJwNcQjYMJYw+M12l3y7ALG
W60iS2zbQx+pj4vAzg4QYbgJeEc+pcOW5oxTM51N2EeOmEfRUOvSo9nmZmlIBqKj
3oIqgZOEAs2ErrGR1z9FbyfFhoUfXbSiT6NuJ4OtcPVuS4oGPo5hx1h5DAw37EHd
PPE2MmmrlqkLMdRxZ1JeeAD0Hcs6bqVmBftojJLNfnxH45pHqsaGGUodkrjwkihv
w2ZFOtDEPM0KIgYl/QrPDYwdkW8cMLRnvNoSPlKIkK/1vok95KoInkjXkUW/y9nO
y5YdBhhlOB0jOMhlJsKadMkLPHjL9Shk92IyJpDaAEdAAvC/cj+UHLWkV0GB2kBy
Amnh/eSjbDhk2yMSylAheAjet2TsnTQx9SDcSm77OvsFcHnzrzJ7A4kTynwl4lH+
/6YMu5sSWmS8DypPJQ3sjPj98pi5oJwRCvKCE9wHDiKGjepb6N2Rb13QFGU2IfT2
yyV5t8i7MCNq89EoODQjshE17cEqYLNlTTCmLj36QIx/F5xYS5C1wd9rA5SE+LRE
N5+0fq0LBYnOEBDLRnpC5mPjjHceOFBIt4OCOEle0PlGfop5BAGXiN2dtiTRFacW
2DEO1Zd0WZdtY+qmm8TnpP0tS7uiFV/skO0VZJaCbR1eg1uoE4SvcfPLJjoFyxyR
v9c/Kq1ICBwVOD1kw+OPWZuVCjo4IKLfMHcdTAOGobkSObKE9SM5botuHDja7+4N
a0MgVcU3Skd83rDard7yRhhD69JPNS4PQY0HlFgAylkqiP9166p79zc3P4KVBSix
sKoIbWmuqgpXZojjxOvLdiHqwg6ka/6/7qG5f09LtnQmMuWhHpHm2Fjf/xvVg+mo
FmDX+tcRk5rSccMA0wucMIdyQWbwjxhLn51RC8Xkul9E//iJ9TqO0KWmwRJB7HgQ
8lOer3L/wvSgA+U6hBrSZsie6lVJO2cSKyFKiZPAiIWvwQpm7y8KVxmNuzVCKuYR
1aoj1o4sjUMA07D3K8G6qYisuRyBYUlu4xhQNMu9OchTHS6GZ4ZAKruW3a7YLK/u
diInYstQPajdxI9C3XrAcqGCLCmnikf2NK+yHV3zCKbYkSWErv9HvghsdRHNAdNF
EqDuMe3ju+aZ2X+V7wT5id9OCwyufl6E/kWXfHbo/bZS16LQImt9GePZnurad5+T
1BultLp/2QktC0mRnOHeTXr2nO9cya5ni0pETFv3bainH0mSpUV5OQO5tk0UCjBJ
pOgewc8jXy0F/qothqhKHnpdRcl1bZF8737hNxIZw1DlYOontSEu1Fv1Agso3q45
cq6V3lj3xfW3qQis3X3IROwr70Qogv7Bvala4Un2Waj8ugUNXVxrCeqoA2Vocrhx
+gjcdGIDEuAdImFCcfR7hLjo3m/f14tknUEeqsIIuU3+IGQqwDOmTnodcF7NFG7d
hR8cnrDPwn6zXr82jFAl4sNmeOX1jXlJEW4WSBgD2WJAqTu62uwD8qDLsVyKBdD4
z/myL8hGt3n/MyXg1G8qeQEJv7z9qp6hz/8Nif2cqtlytMq5UDENpA8pUjVrZJIZ
UbzCx5CWKFbvL7bb4Svsb2CRntG6AxD1E+ExaVfiO/BAvYlzrS87dW2GFhNd9JQM
MN9FkbQ1HI9498YW7aRlnor1ST2nRYdBt1rMSkwNiSUvsjSqXLoxX0/kchgYjMpw
Ehgdw/K7eHtoDXfZNbpLYBL3GXidrp84QkEIZNFzBtw6WlrO9/wk8DUcda1ht6wr
ZVwZMKxSxUFYitus2ADrAhMaeNeO77UY+pVprRE34i3wXjaAycdLhWi3JVLzA+q1
rm3ENbtxAW/78AAstiSzFZtj+22Su2TWfqxI1RzoIyl20lRnnTIbbrk/iPm3pgRb
4TXEg0DN7M47LarX6MBLTVJeo3Z7GBTUe/INA9Mt4SjI+7R9GlurAPW1F3aOvGSL
Lt8V6k87/Khy6gJTraCrkKNYp0kFXz+CcL7GcqBuy87NXUqBxCjhSDLj+TjuzKdC
GpgZDOPfx6VtKpWjdVbdjeS1VSzpWeLZgwPDuLSbJ7Pxkuyp476bWdsPxVXeimlp
J/oOjbLtO2v6Z2b40RZYpfOZNcPkGHhcId/oa0pZ55maXibk/k2t19bfynHmxMPI
5SYylvdro6ARymxswuKrIG5f0HRuIAyi0tj6m41+kDSd/+Bt6p5rlVrgQoyrT+PV
mFwni3smfRKo13fAw6QALK9me6NmwEN+f1N0/nFRikV/LTShq2vjuX/0xRVSCwdr
NLahQCX3sisLSMaFM0pFlrscK7gpWr74rwM3a47WkGSU+98CVQMzdaGBdaMZOc9R
A/Khv2BjpUjcYbmg+nI6Fl2utAC0fX8Bgw4uT5Ib3ZFjpb+CHTUzlkA3bDmrw6UK
xAxNN/fEGOSfHw7ywNzHJxZ9KYzrfyrmm14ewefU9v1UpzOgvlM2ZYjIIZdDQaCx
LshmQdN2pUJrRh3H3iJgfFX+GfnBQ7ZVf5lqKytI7xszjZZMllKiiXa+9rV8LuLY
Oqi5VRWBLnkQ51/YSLhJIuRSEHPjZY+8zmamMGuvYAgwtTCc2nTz9tIaj4KoVGbK
Dw0086DVHx0gl4RLLIYBNGCpc12r8Y84AaCpTxvHzXdNr60zsKHsB5aoiibzwsYS
kRS1AyHejM0qI4F3aMWu/YB/ik27jONANphq2zumNwW/r4Iw+qYTnY0R8/inA4G4
uZlh4j+/wCxFYaJOTQza1RMA5kL5jRDPg3E+LnVmiGcHQVRCtJxQCCt0rMl4Q7Lh
phGWylRWV6603IV8b+hJZIFf6fZL4HenkLaf572syi6G8Xuf+myo4Z8ztmWLTsQ/
vZHjoSY13Zwlluw0sKQ+O2AtTH3/QNNi1Gg+71czhoiUlyt4PAXy+SatiIaTV+L0
xD7FgDEXffKsMLMxMnOxtuTqwo8BHneXvc578zJWDb+exTfVco1B4PUJalXLlIve
INJ2OKvxYVjXijQDvTm2wEVjjL4BY3rBpMkGh4C1eKiILRe2SnAjvW/BiZqKpCpf
o/IbpCDXfR2OMiprvi7o6oUqtWgUvrSQ7GoJKSVy3F25G5aNSusJSoWjUt0lpzNK
q/PkDE7Gj55tunfSKchEj+nGZ53C5Jj/FWD86nok7fMUQxHvIKBMvji74/FdwEfk
UCYufuLJu4Eh3/y/IHKbFrP1x4p4ElNx3WWMssDGCs8P5BVQ1Vl6JxXKuduvYUIl
RX9dzuCnEQUDiu3R7ydSQgNyVliD+YvPbStl9lihS0OcycMM+ADTyXAtc/QvWfQI
5An9N6LufL7x9/HBPfd8hfqgyW2v8pED8wAAcQjmsQCDRwB79qR6yUefvvMoNZm1
Jb+9+jVEKg78692//S8e2LpuvJRlRBZv3pP3N5JWDU1/ikHY/r4eGYAn5t5cIhuE
0A4dPxJwPbPcfzdto9vfMM0Ts0asQjrMZLy5QNdw+05ldhhhdgjPo/qiaoRqbaaC
cA3m082p++SxeUbggmziJ/iqdR1Hd9sd1DBsxxqAztYRBw9koqjmd258pHh5eJkg
jARBu2pIe0Lqg5mk37Z2XJdhyl2ayp10fLJafN6HmvZl4YRZsvSQSQKnLTiN5J8o
+MpdAcBMmbdKqxVZpiwP+YndkZSDBtntBCR/ZFvkSyWjQwLNGtJgW7JM58HPYQCJ
GvjfSB70yPGAF/y/zLawkwrcZ63jjkTFiFH5bgnwKny1Mvad/XX1Vxkq8q6Honjv
pxk0ya2VnRyNSZCZRyAe2rH/YDhFYdSD5yLRQjGLq1T5MxVcJ3coTm2FS6ciiEBT
GwlKiTABVdPqmatQdQZuRaKk7A2kYzQ0n4RKPbhP2hY+YGK1VkqVsoVBQP8ZS8hz
HBYKWnp8UZ1ifAp23H5FtPk2YBJO2M5zRjZmVIPnWW8PX1CimjTjIoRGdmyYynb5
BXLdSiGLZnmGw0NIRdhHI1skICrgNvcqVDo1NaOBw/Qowzr/PZhdndlvvPnE3IjF
i1pfRNUWBJjEqZVyITB+O7YB/MBuJp0RuSsG/8MzLLhd2cpXwT2UF7qJVh1baZpY
RJ4nwSFW/QJyJqpsb/g+o9TCKcfcdyefwhDFm6nhrDO8FZEqtJGpFZS8BSX1sYYx
9wJ2g7GKnkp8VNnM2HVVH63nlzqY9rlum4uT+iHZ1j4ICpqS0WSkOOhTH6tRlCLA
JtA3NGyyRzTiEen9Sz/1v/WhCTfPlwXszQStfH8Mr+axSeqT9JR04NU+vNtG/T0i
E8lPJz0csU/w4brCbcn/6omiBv8O1o+DLpCPED9eLnmNY9PH50pcwsdnI86xNJq2
7BW8SpXDEpxH7uPaf38uWnAYC8TUrQQFG9Yj//5rrBS3gNDOFiJ+mIxpWoXQb0Nv
7ftLlLCHB9h4aw5BLkUlFZECf5QGG7ZqvSYdk41GC7TtvYOejGgnJeqMshg4AhC1
uYlqep1OtNb01od3k1trN9BEe3ROCzpLa8ZU6NoFWj0uQ4+nSbChRfyVvtmAI3/3
qsgtKZNnmIXh6JnqrpeNm4TJ8VvCB3h+xZzsNMnR13+GyhtloLQ0YElvh7P5+AZ5
KqJPq9q4jJgZhmkl9BDhF4mw4cAu+4UQXZTZrK2lheLH5lePP8/VsvZtB47yu2L6
W4p2X93JffIS4QfW8555LASb6FAQD+DOWIHWUzLPP8umJRk8sPnuK7DI8+qhtcKu
7ES5cFT8+shMXSDDJlfw/4taEI41qxaskD5unbgxV7i1KyOyYWPUqfbs0Pw26XMM
VFqOqJRtJOKIsg7a0Dj1sxTeZCYxejS2z1hnV0ixP7K5dB6moFC5AYAhYOF8kP+g
x/wUZP/t+xCwSsYM3gaF2SwDzBnavrElEnSSM1GgQCPQIXNyqMig1OYB0I1djplQ
+emes8hb2NeBml2lfm0z6kY1qKsBAaS7Q+7EuNRf5v1H8+hpYhNnS5z4xGNNfLDs
wdyrfg2Y5V/yjGbGKcRJ3TbAE4yngvvEPNuYkSGOGwvvdW9jNgNDQAqKeCaxXU8P
prr0w6aNkjy7xdcshvmzxjnkF4xndzq6DQEi4Jjn7W++7wOyeeVOkOuRmUTLI2tR
6lT9FYFL4qkDqdgHQp9nBsyJ0Nbod8mhx1WkoCwn4HU6DoTcBSEa737ER4eL6n43
Ng0B/NWPh6rb6VVX5b0WvHkbCBORtvLvMxzS/OC9TLE2ov8XBeX+aISP4a0rSPwB
ghffzbSg/UU+yukBGlerQaHd9CzLjG4E9DXYe6NlLO+AQu9BMTM7TAJULIsDfmD4
jQQiqCFjgoiu2VZH0ZGp/UcSAtwab+naRHJohjZI0q1UbmPVE6+b+CnWbdkdggmE
E/eheifpvHW+BQ6VSQ1wXlKDP3hEAhOAW0gZyRAhedXXnpHAtjpTtqjenE07cNBW
a8874gP/xodj96fW0StMj5c7XaoTfXP02aAJtzaKJaXSAK7MpwU53AsHkcvj/+JA
Q+p7Y08+h6vtjkKBNCV2lija/R/EfdI+3o3eG1dxYfNyeWFfWhUD9rKeDzOPzL8N
bychHXpRmmwCEvQu+LnsoXtypIaWoAeCcyYUI01Kcs6g539rOoJg7kaLJ72ScTce
8WXVbEYPFRj8/5jYrULFuDMAS3IIAZiSTRBIlf9FTCLew7XT9OgzBa3IwLUbFrDH
HJzeWCG7sorcJYqHvW7Po68OZD0RVeqTfRRK59DzkutBIbdyyDs9IqeHyAW1hYEt
A71ly9iTKGtiTUfXBCB6IMVUc+VSea5mI3shI+fBwRpEJ//1qAXcsOsjzjmH3ctC
RnjVv348T1NJ9Qcr/sT1sqEx0fgyaX73SbbMWRiaZfQh0kAq5DmtMQffR/L4hwBG
Y+msjULbPGvr4v2I9nK5q0hi59D7kbtRhWR1oAJsQgbIrl4QaO55h6D9TdZXPfoC
BWtzoS4lzhJ57SRHpj9rRchM7uEPqy0Pz2qOfBHSPvQ8yuX1e2nUKrchiCIvz7ra
tydCUaFFCddS8QLZN5iqeg4aZWeGUS8m86DRYofkkiF/IZs90XxgYNvJjLwGHqE5
TzOlYazF830YWe/WwCTCifYuMV+jm1p6+EWJXYPMy/tXyevkCk8xRo7OGVVVCY0J
zhyJuxrJWgf3oEAV1bP+7PZQ68IwlEcUaHCD90rJVdnh6f3N+qlTibn3gsRZyg2Z
FeNYmIWBplt8QPY5IEjklQfCH+Cv4k+xM71lMZ++qajKdBQHQil2vfhEt682RCYV
1AgsiNlepewu3kpOKJruJhbTa3vyCZPVEIXGqMb93O9OiTZLClQieu7Oyg5n4JEI
3PvtiWwt6oLuRjC5dPNuTndmFTqHj2ha07tbV2AR8bR9GbfDVuta8noLL8a0KlYU
5l1E5bPAAHxsHKZlaniF/GI5/0GvybmpqMYbfU0rxwue6RLcw0PsSOt2P/q7nabx
LCF4B0ixeXyB5/cs/vltYkXsg3Z7PnVS8h15Q8F+pILgTTJAxrkUg+j72Ml0C/lp
JpvkG9KZrKdm66DkICEG/idnoSpnLpU3i1NzKdJ4PdsthLNO3NxRJbbax29V44co
9/QJBWEcA8oOXhIFKX2699BM+ra6ydlKKM3/1OFXW9zSJyrShoBUwWcSBGBDJT+y
3SsBmv1UvtdrBou1o6Gzs8UPfK97e7LCffC2djc4Rv0ENn3Ns+ukCl1REzJg2Omo
5LLmTcVy/AZ9ef/pJJFu0ddGzZ0s83T41cPP8o6VKj11XhdabzV8pHFUdgP+5X9c
kY/KdExfluOv2iEU4pbse2zo+ZatgA+gRUbngLASCYKoo6RF4UHlYie/CiPCZUom
C94NXXPR2lcwGHBK08Xv/PWU80B80pCJP64mYgFJ7tR+f1iYssVdG1sIvVylm3I9
XVa+GOZ4ZTmYYt3in8A0ezxpJ6M0ep73/l6ue8TDxf1G+KfPmxBvYUwZvAXa84ZW
RRXW8NkGwefIGwPAi0e19L9xNoNUFy0WyXoGbogZvT1UhhZBUsbXpgEYwKIZkd4P
kRwCOP9Dwu6Kobh2EbNbd/3MF4xWnWse+AB1FzwQVlizXwzMM5EGMR+lX/rI6Nxg
r5INLmYX/z4cqlET3rkgog00/mrqL5ZC24X2i0pxBdksUx/y64gob+Rk+8aryjLC
jJkqKYEAfQUDq/uxuJg9uknOgkvQgmFjefpbE5CAtv/YyvHjs0YyvHe5hzege7TB
JzB/s5lVA2KMJc8oHVkXv95M8UHW+3def2LD3Z7QcKwkIJz9sAG3+/6fRyEW7M2d
pMK0jkUwyoe3SLKc8dAH9U24XhYuDqUr8KsKnXHLy0gEsA/pW4vd6BqZ53ymNGB4
OjRXrRbLeteEXa8y+FumDXu5FtfNvt2GjzZwE7MlYobndqHJ3DX2ZeeBrIIUd5aX
sxtcygPzrbOpyMbpfISt6Dts6QRKWKqG557cpmhMtEZvbCR/4I/kvUCg2K0mRH3e
UBdJqDyiR5WUuyMIuDM3rOhEz/he+3WWR9Z923gWGIDAbO78eABGi5yqxbjQMiCb
VYOZojHaIYWSFSsw0muUdQTkLFL01oXFNSqcslulLEg=
`pragma protect end_protected
