// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lws0MsvEbEe/5AAXL70Wv8xKNyDrpGmqRcRiq9LTBvmT9bTPT3CDwzZFJIxseWUY
8rbs5ol7fioWiACrCgf7L7fG0HnAOZFqZwyvuZofZY/3IfFoxtqXJNtdD1Q9ZEJV
B4IyILWqNAP2SRTEnWp/7SgWxtbBjZRsubbZQzYZlTU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15504)
XhkOMnncLAlD2zYieVWd8q1FlQkoUeOMXeyCSoencBXbTYmhLLF/brSEDnd4tPc4
Hv7g0ShQT8O9VEZG54UxoZRU5HcYWO0ph7lzRdB/Vsmn5P/0xI0D88iqS/QPSsEV
Y/rPHdsZ4/qm/oESKyzo4Ha4tn6QUqbxwAJppJKIU84m1mEf7V5t6lVU86ibRAcd
EeYiG8q+IDHmWSNgics67yCFQHPVNZZlvb82OxTZty8SSaxU90oRxNrdQQdkquAF
cdTMLoobSR3aXpwDQN2IvgEA0zY4Pcx7ob4UsnmaNG9lCX/iincELSePk+EfYL8f
jTu3qtgZIVIQjUdddsiBMUeroqWoExNzwheZP8PZXoy0LeqWnoE39hGlQQ+7MnZR
w3RY4lcnpZAObx/rdEN/TthMGSbjGEmDrEIs8D2m+g+S1vHb83BrFC07RO6XDvXD
Q5FQEZalxRMvxtNG5j3XsbzFk8A+E41Z9hN8rhuzt5L5OOxKGLRwBiS6NOgPeMvc
6jtaqSXT02OQCzdsKgLFyVEOLIJh+Btx/OAgqRrqX4J1nyxKRdKfRQ75ltZeesD6
xp8c2V3srLvgh9DGgkjS1TDZe0ie5iOUTzmwM4n31D5nN23eCz59r9jE+GKmj9s5
qvNF9Wdxrm7R5oQrjbsuDDXOA2xFQ1OhVbhs3nknTr7Sz4dSbilV5+AIXcUermta
HVD0m8LHxFhJ4r/yaFj1YhY9/9JHGQ3z1vKoG+tBV5LUC/Sg8z93J/ulIl5zAx/l
Djf0yFbt28/IIfEKpDxX6aShNQzqLYFIcsAq1uNJrxpMx4YVqNMWZ8m2bMkb2ged
tp4RaEN9ns58R5BtFs+ZYaeFtWg/P1dCEnepJhS1JOVnGx0vTdzUqI3abbJ3+IjD
P6cvmctctk/CoXNWR9oc+n2b5taIDr60wQ4WOXW5sgtywvjxGR5j2xrCXmwv7uBY
Pa6tmyBLAePPwCmhiKDsYGwBGrAynHB7Ar9JZojI2zU2ML1E3bohA5Pee9Z9EUEL
ktdsqm9HJ4D0sDmeMDl8U7wE0jEYW97P0+u8uNBgS/yOcHy/bEp3w2Uj52cU6Ybz
Z8mLGCF8FneoSx3nOUdIB7DvX7l3JXHD0J/q8tXgVmV53Fj4wOC5sn8g93BcQvyk
86kUA/a+/PDIPrhqjcGm6e/Mx/0oB6w0tHD5eatoNLpBbS3Oh1O9UCxTm8UK469G
/dQagfnVtBcd5vdJ6bwkkFZq9Ib2bLYVcXS5JmQiC4zwO/MgW66QbXYINK+I484p
2ijcBS7yVa6cfoenyQz+0CnMNsZ6AlM7SPXbKgJCw4JJfPZ4XH9DKx7fHskGd4MR
5N4QUB9Drk56VXnZ76/whlW4ifTMMjzYbII1xR2NwU3zkVCl/tq2N6P9jO8/sdrA
WGNKH1Bwv0Yc/VyGVX2cq3kMIjeOs/Ec/8XqegeMFptG9IAD8rNZrud8d71SSBo+
V2ZU7stOKB0gfUSanHTQfMOYhsPb83X/xrJJUtRdRe9/5/t15JV/TxQLgnmNSrtX
rUzLm0mqirvgF7G9+YIbj4n4R5tqONclTVppDd6CZwaGVFtTBQ7qWj35icX7xwN0
dpbKRUMw4jqcnbN9eP7Q8k7FGB5tErjAMVpQscNMyNrUuSp7CPHRjcezoI4GH/mW
jMPEYgYyK1MzoG8lYt9myxYUsceVFQSYoMoujGlRupdCbzNFW972Q3A3bRHDI98B
CusOrOQsMpxDTzrDkl5dQe8qKBn4rJSUh38sVpwWBGSsUREl3lMT2304qb0Twwac
+VEsosJe3Hqap3PgEGouIt9qc7EdcJZ106zzPQDqi1jvBs45e8CDuRBKPez+M2pA
ImklshQXDpO9G79XAQLlaQi0C0GBCRo6tq0ehFRpOmRbFB+TfafHUwtSQznF5kJK
lkXGsOXF8k+b2lfEu5zZ99nBd88sdbP9pEUYmrO35JlTilFltQrgYS2pRY/bB/LX
eU1sCZ1PRwZMNQJ0Gl3LKvH6u/q3WKXWuYYyDU1ma6HDAS6mPnmGlMZYVIoTbk8p
wUFvWeAsnqVvZyulr0bImdmbxBBWCwRiTQ8ZIs7HxKvh5IFC1Ns8ranICw/sfEn2
RbTq/+o3TIomQQQVBOu62nKGnChbULyABXj5zX1Tm+JM4tO+yTxB+UCZ7n58vFNG
kr8JLc6F/P3NnZ3sS7zSPsxr0m8ooezH9Rr9dNvAR4DJ40Rg9Wj40N98q3eGL4F9
f88za2IyMuvFTPnUB1bSfy6szBLKmItl1pJOR8xbuo32UFQt/mLeR9h9i+23Bxxu
L51VFqXPs3N3Tf5oM10BpLpcceQAN2xVJ56HIANrOwK5Xses+P2V8QZDjVHOLUHA
pJxdqA0DhcEc7IzfIUdRjjY9PTOhgid5B35IPh3OLAdsFgvqxuX+JZp4Nv70eS2O
dGRDmUDf+MFPFUx6b4E3P6dj3CjtC54iU6hMU0AGmDYguWnh1HetgqcAUNFxPJk2
8frhgHff+TplX6f4s9Nqkb2L6+qGV8IyLCumfeQneNiktgdj6YtjoH6/aUA2zno0
GRVvk9VkSckckv3Y5ACqTM+7THNjmPcJ0P59xzPk4+o1IcJA94T5kCGNnYhO9wtt
clX+7yjPrV34csVjzil1lsJ4YGYX+jEjZvkQAc83ry9c8AeiILeHSQhjWgwef8cH
ctHzdXha7Xj6Xl9cSPeF9wUItfWhLyu8jVfGzzTkBWylNGVhsboSyUQ4N2K4sFJg
Fx5n368lB0nqURZMfxGBu/m/1xxOfH6NL5yhhPsDq5VUFKDu8JLiZWt8JY7fxEq7
zgGSypBxqLNhAWB67/0WNUspIH5kSnc5cDZ0NmOMXFDtKKKdET20180uNbn78w6H
QUTG3OJ84JNPDUBxyFQXHyNxm7GKt7P1/6NWfU2/x+F/+P9lR8yBGv/3BLoOgoVf
G6qgTjwkagySPgYz/oSQM5g6pmXZ8bJCZ2TxMBuwZTzwIYoxTBXg9u6t6r+8YgwZ
tzNxD0BTo9dqH3QdSZsc79Jq/cTEEbI1DcqKeeLy3+YIv6Gn2ExaQjygvQjVWB9D
HC8xbF5dYKVoApnGy87su5Bw4fCbvwMIt0/gtZ/DlDdm9domFElPUGaP9v5BX/NS
kDpnARzcrOOs4fcxkFSwqR4l2gq3unKsFs1ftdvD+5NPc9NfhDKDdaqFsE11UReA
pxcxyEOU4j81eOHlRSJxYfYebfaPeprQxIVzQNQkodWHq5rPmJG8mlFQsyh7Qgtc
V56c1Cz3+aiL6Rv7CwkunQ5aUH+Fqy0cDY0iyXEL5JA7zp/77p211SqQc0Vs0iR4
8aDejvycj2OAO/rL0iIR/zhpMCdIKBnthG5cOksbpsvXSR7UeRFM40v5N+nzS7Dm
2QAX95EIOvDT8SkqdhiYGJIj6CifTcAfk9PN87FweeK+rNdfOaMbG/K6aZftkSew
NgvMg7tbZGRqXtMGAEsaxwBHpibGko3CJQXEJtjoRuiACKjKjC+QqqAs3Gg69WVb
V9f1ftQqNyQTD0SbMy7S//3wcW8mSdvr9mw2EM+npWtzqO6Q8D5EuEGrZGGKTWz1
dAgGUsvfT1lIg1e9f8GcW8UQP8kxVT0gnKaHWErxvBZw51dOUaG6KJgbIgKhRN/p
I3MYCermLnmcV/WBIsfojHO8wvehSmk8XMWf93cl2l/sHn7n+dQWOBgZ6Oq0B5fB
TbPdIO9k3Qd8Fmf9nIMDV6fQIuac8FJpH4R86VI27VmYv4cirttjYqhyFT74t3qD
e+kvmhEROJ3MnpFHHrYTHK5eA31vhYHrL2Cp+2ys4tVaPUI24NuS3ObiL82zpK9K
bzvt7weCKP2m0ZtDx2gOja5OZp2PPSza18sddGunG6b56Sot+gTo3Df6VhRD/5GG
emXWnnmGQ5Dzk0DvWjJBxyAtI3Pey+fqQCu/3ztRPYEB8lL9SOenMTKnmQRq9Sgv
B6EZ9K0pNWnzNMlTMJbBQCn4vI4LEHBcMp2TFYFeJdYBe2e0gQz5PIIBvEGkHA77
hhgtO4FuX5ZXjCTt3VOv4RKhoiGKkUvLbxN4RlUzME5QhxsmbF3HF1eZSI/VEGP1
b+ie3mrKRTAgp+C4IxXmgRGFNRAx5K8Db1OmHKpa+HO+PTHNftV0uiW4LkfXnMlt
/IIRST7kQa2YAUDO3i1OVjc9hpXDUtKlZ69n9eTCOmIgkdd5FAqiiXgR87OiBtsv
Q08H5ToawWTm+QoANZV008uzT7QfaTpBSgydb/uDr8kL9MrAAMZCX2PjZ1/bMQOa
HQG/ko0KuhnLeBs4tOChZ5FU7pqJpOWpjNebYqTaR+qQimiQWStyvvIXE2wVIqp5
690O2sFNjBKgBbkw3C86JVvpQLCUyNkcBISnKbx0ifNVnrEDD3m38XRiK/UWVJjn
ohZfhFijsc55ItdTOIiepiYunZK7m+DW0eF3YLdrnqOhWIEbXJq0cmOloWYfMLc/
muQ+/zNQ/JQrYRtLagh14QpSy1+gQ2ROtrcgk0HOG+DeoOIg3X5yjq87nEm8nIY+
CvQxenLTXM77kgEoQn7UmTrGkC/GQ9SWhn+7o5uYAy1hQ5Uhplc+s89Fi10/zvpQ
9wBkKHlit6uA1kGysK1+Ua57geZgsKQTx7UUpAxxyIE+w4g3ai05uZqdTZrus1BP
NHxJ2Iw65axJzkTH65uhYjt+33jfs+8jYlswgPz8vEgupiEvSPkJ3ehFcXIO71n2
URowOFotWvQJi1bt+CSwaF55XrSd8Fuf/oajZ/9MV2HqUEOxggg0UIuTcHLiTcG5
zFinBcgGP44Z4LhMJr5c6V8pCLzqFBu4xKzitZMSOdmxezhcy9WSi6yDYXN5R8QJ
PBI9dnHX0z8pqw/I634GWogPvfM5JaSUht4+zP7AiEH9hLJHpqRjGcCkJW0kOAy+
WxR0YsDd1SGrrxFKKRvIo2h2AQ59Yt7HX3c3Lj4H/tnKPrivAGjM7FhukEr50sOr
EdzPgJkn4EsHIXeLFVb9qnTxXmDAZC1vryrslnNklaXyl5I1LqAPo3Gp5WTNiYFp
TXO2VMQDSbG4ZVF2+0uuZ/cf7q0A6wHOZjExNhv9Q0WjmC3dkshBechjmQFIorA7
vjAZmGu2R8Qi7hDqMH86KJKtcg3qckOHC8xHaNru/04MU7L/CyOk2vDboVOX+Yvz
3O1Rm9kdEPrfuKlG+f/0HDtJ91kk5zuZ+mC0jGVgbHCoGfFNlw9oTKPtmIS3a30G
ZlJSJNm5xPoi9KGHMxFRYtkVkcYhxcY56/RK/7zqBlirXieKUS+KLrASdLHX+XsX
aWkJ9YYQ7RyuQ1WhgKrJZPoe8LkPkDFVdQtXB/1Efz6CfwlLckhtVkFTpmKnItxt
VvDB+7OYziOz0Xqlpe7rIInoOHVNBuLaXkvIVLYus+RK+vNATSh3wGoffN6uncPz
ruo923a3jd0Co+CQ6vmT4otE4FXBYm6QKyH5HoyHlVchDkxr1rpWkT6LRhxaKbbu
8x5p+kEOv99uFEvPR7KkWf5qHGDgZqg2/fEyb4Cfp6tElK/6Yx/a5VDbmyDUlwgJ
Th/321SdK0QYOaPNXN8VBESJISemYwcfxAwpf4CM/eGMSEW4JAx+viZusqEjW7Yd
RF69c0z54XXssXpSLJxM1fexEIpacdDYZvLsFsstNUXs3KPMy4G/mxwoQCrmVi0y
4C9oOnhuEl8OnM1G5rNgq0xFygUJIyIWdsJXxxVOFq9vS2hiN1fvgQKDw1aRJGcv
/XDaRoaYZdHkoMfecvU+BrUAI+nwlMlHFPEx5lsZDNrjXwgvmkrdDq4y+ELHnHn6
PPr3GdKDxFYlje78FjlC5MkPPeWxm6d3NNFMhiBOoUuwcrJGfkGJze+909biXP0f
HwDVFwVWVVtcPa8BCS3OTb4etmPW+4Pd2ZPet2ptzPF/pFyhXtcTvPvyWDdyCDG7
1ALL16Fo+6z5osqrxk7mHvJuwwH59bWmRIuZHt1n3A1DaVQsCzami7+H3YIlj562
OM0jG2azAKELiKnBRIDXAFTdHunzqOxSdMc651Q/TsTaBDKB7d5xfc0rQuCZjGkZ
ZgDnEeuuBqVJSPVbulCB9dNU3PGQjiK8bjd3x4iJ/Wa3iDdl+GxmLzNN9y1hwZ7r
h2clav/YJGwAsHBuoriOLKOcKjR9GCYoUY20Q3AKLcEt+pgTmmr+Ya6tDGLaW1Y/
0UobIgJ3bDwwpI+OFHVIN1Fq0RAKNaJpOkdtyHOfsYt/p/7eVG1ibxpdlal22shh
/KWq2p+AmbaCEJpPr5qNEL2LryfZUaCSjJAJWdpAq3U8FIOQbmsKY/V1oZqFT9/I
7oLe6MRx5/8udvv+Wy2swKOLPss1n7dmJFXOtGd8C9pWAGRSqBhV0tcc+uCu9ryn
/EMB8XcEJ47ZUZAKUKfvt8M4oh98CqqwQWdktYlmvSdNRb2uuuEJwlHcTOHGOW22
hZcWq+aPOZN/xwjdjJTPOlJvUU/DKJ2ou8jAqetC0vQfG6E47e3XGtQPTSdQ/yrK
9VegOMUBjnHYl6aIK87tHWvR5s+IabPNir4bNI0N5+7U5KeT4W8GyS1UeUys5WN0
0RFqZHH8b/ufSjh1rwtJgcsiQ/7cuKlZvDxFZpIjbYFkSzLK0oNZxJPCHKJWKQTQ
S11IPzmLFdSWOjmZ2Kgbd5mSP4gst42oGtRculG92EgSfTZKTmMsN1t2QiZo15N/
OafjGanpWSb5kvxyunm4XbEBsGGR0RuCpWdEWGEaFQ7TFNgE5f1naFuaj+wzQZ/h
Lu2K8tFmddS+Hmu7a8rtSzm71c5H+ozGYOJPWoh2g4GNRhn+tqBUQUzl5AjrPCyP
+BD8bNM6ld/dihrHhrfQl/YxsVOev24iLffaK8BqaVu48aTM8SQ7qeUkAMaoR/FA
vsE3buvrKkgzo6JzVkIlHbVbyPTYgBbRydOeVEPLvLACaDDb78kN7S0rBXiNpHHQ
J1lm4Du7YM/XYbIFK7GcrajfeigzqjhfMW5l7mYrgi9M0SvVeaVn1eCl7SUz5x7r
JtuezDr0uN37EC08Y+GeLDFnQVSXYsVsuAWtq3wly3tPAd/tDNb9CYdIzLRGpLZY
pCVgOjCyUbuuxOCKJoypOSG/Bh+KUsFFhxsgJ/chLTNi3Tv8frFsU1m5xhzwaWsT
TU3bsdugysHjcea1esDIDlFVPqhFTjqpjp94IaaZQaaQAWTeAWNFyUXhoGoNhOk7
cSe/RazedF6TQ2OF5nijQgNS5x9cZkIJNmNODJdTSX3QZBmbidVhf3aQpj8vWLjy
Jehgdh+PUWCPHTqRaTZKqhjlCLNm7eZSr2kV5tp8mFn7+Mk6FRGN+uh5a/kMigJ3
a4LNdocJPMR2JYeTWqhrZPn2VYZ50aFwMOW5Bw/hQMQozd1GQaIU/331zodQMSin
M5mkAwdQXfy8TzpoRQE00vEcCfVHLJDoOZvi9TD7lNtoshTMveXf6v/iY0tK6aw3
Ft5oLZ9SdYb3vDHmR5VWOKHoMEIe1DjqZbl2e+GEw57qhAoncPpZ0HBpA76Z5yV7
a/++9oTyxXdNy7vxvAmRpJAFbztwSMvwWRaXko9xZzTNA2HGFqz7Gn/pme0bxGLm
j7oae5V27CWDGp1o7faDZ70O1K1faQV2Ldv5idyunQGzRgjZBrnqTcu8Kym51sbQ
T+DpSScZoUOJ1X0Zkpxg7Dkd9SLM7WE4Cy1H35bkAMNpSmfms8dCW3Q/aVnlCD+P
Mo6TqBn9ikL/M4ez3q249Q9TEtjOn5khltLVA1EW3FtLETbkUapfF4wGtp4h27ZW
KzwvarQhwM0S+XjxheDzoXNipDey52c7GmOTJeuHYKlVatiwx95GFka1lecOgtjN
+jvmXwhuHTBc3s7OwhdReMw/XSF5+Onm1c1BsRPM0ITVayaXh6AvBxV36qZM9MzT
H+onaHeTjOPMCpZBeIuIGJ+21f+cQAsA35R177gsPHpXAaRg0Xk6TS2lil2kG2vQ
thGA6PwQOvUThJH6WrxSfnHNMugC2UNdJeu7mrSgdjFl8BuAt8rKTRxQU8Tr0aRa
HuY4yqLegscg2sRrDHEw+SWCdXhCuj8fVYhouXm9lnhpRT9mssgUdplr4SZvoIfd
TUjcTazRnNwRjbyM/FcyjE718Eibock8bLOKMV/w7oJBiWTHIFFIo20xv1F4OMpo
pF46jH7Q2Dol+J1YnX1pVONfF9d7xwtOSXktzo34nqcyzUhQsT+ht9PTWmDiFZX1
x49FyNYE1sjV+0sGNvykF9e7oV228LYZzLNcm4Iwn6js0mPIobd4i8X5wtP/yo/W
wlYWaNjib9zngqwqDedntO6HkzFs8WPsY/oaqzGfMUSSa5o0RzUhN5TbJWdpOtul
jyFcs2knyZhCIcAnR9FYuRPE2s5dSE0vSvTAahSOB6Klcd/CgMaHYo+lt1sOjOR0
85fMEaeoKFfO7+RxYtVoPFQjzQuU7YF+7rG2VsuM6UKdYUMvS6APQ5tyyUXrxfst
Ujp3Phg/UbvCaki4w0Ya6iS8WY/AKHW9gT8FQIgYQOHZkP+uFuMbSN+WgPEoxuHx
uwiA5YOnnK0jF7uUSHyQ0ctyh7805KmBCpzSx8P0G8Djox1W3liUPYJv35GECaVR
L7O0gjSMvz0ZFn19n42a/hx8ksJ+vhWRhgs/PBBwSmGJkTEYiPcKermIgK6Yw4PU
P1tchqUPmErkuuR3tYY/swJTqd2HZaXfI/W78M8fUj7d2yFKqmuyN/JHYFHRzstF
D3Hi6fXQRKnlT2IMU9/bM3gzcyfWWYWGGR8VKadAK5vUthX2gqSpPniLY1o1kC9z
q1UMkLJyJ5F+6PfElfodOiegYmQCENXnEWJmqA+gW9G5bFxufDuBXl+PkzEKiknL
Q4vZX32XIPTXV6vskIBC81GmCmLaIQ4v56zpi1YN96n1azcrnlbPe1UaU2OeoqTd
MOCXx65fyB4jHYhDA4s3vCNjwYXkrrkkTdxKtP8pTb5YqdLg5o/ijp6/TjzVjmXJ
R+pr/cJ1CaOQuNm15f/hxNWpt3t4PBtwMIpcQLmVrUBjWnR8vlt75x4SpMAiQ9G/
vBewtCe5Psk07dEd5LFI2700WNDLFGfv0/TVuC4U5e9r7g/NLg/hJJ+svgmXUOc8
54KqNv41b/ZKBbrH2bLWzHRGTZ/1JgDYhljwo3aYBx+uMlEhoWpFvkOGu3B/GI/z
JTH8NijugXJPXty92AD/FezVGiiWOCpNfn5izS8nov3QEscsT+qpvp0l/yTLjU9c
axFT2uvsPhVD4FkJXCWi9FdXpKUzej3l3BE4UQR8tFjil03eTaHbCQLyxU4BZxMb
OUjBTxEHA4ieOM//FJ2wfwpYV6ZihVomNmaf3djINcGgSiXaMrylnYbSRgmdSYFg
Y8iRd9ZWa8JAiXRGRqHaO1DzsQSQeXln9VQJvgH/UMxzCv9eD5T9TSwGdj9JooH7
cAlOZyL8PFwhiZlEf9MKFW9XGDKTkdrLIj+dYeCkoLY2hGhjaiwBj8JwMdXyFAv6
KeUVfJWgIfcC1jP/YnJlwoKuZ+TBm1P2K0UtCp7ewgreIyiJPylkeVHYgF5XgO8T
MllfXLtzptkRAW2OXXjxZMk0EhNt9cKPyaJgoRRcLWRE+xhbZu3BkjQGk6SyykG/
FYS/+52zkFLRczkliEfZPqoA4gYUE8VNNUEIh6gYQ/zdfxzdKtrlHC3FfeK4aEKD
ln7Fh+QQOanuu63Br2lFnuRr2hE74Rv/7LHODT1698DM2zC7bngr3M0gIpjXmLtF
v0WeBSiKVlWHLAe+FU+1o5TYuzxVNiD4AJloykT1a2fDJVyRKQfqNMcGMhX3Coj4
eBEOzKU4zBDK7s0Y5GHOYC+jqGmW38v+oM0Ssv4pP+JPLNeSA8GoUzOxNxhI8TgJ
wlg2ZrbKR+3iHzu6wOkODprh8z7Qf+A9IzrEPrV3zsYS3lPM3RTyepeosf6kKbML
LdiHVI2glKB6G0FKWpPqWVGt0Zk9Xu4XS/t3PZMKooIetc+J5qEmxA2BM88qlDHh
fEZtS9qka/y0hk0I4PskIhzTgWzoxirIDnJ4qINbQammFrB1twoIngfMpGQE77rJ
gqgC/9uO/YZAXkc+mRDjABcY0Q6VE303v6IEBOpiOHB9xfL6yFpVJ1tD3drZb+F2
Ddp/utobCWQbrR+HcBd7ka7FFYPD+8FijqR+U5a5nxlymZ0OCsnuPkHNMEL/7kSa
aUdH7hHD31EkHCRbpdFQzhIZAORpl2eUpoDxEpGyO42BZgErZ9RPyJSUjftaafbK
2sDzApz2b12dxupJRyVs6L2BFxmgGsDdZphk9hj0r1qDhLaeEqLjF/uUnJoJc6bZ
/IAY+H1aMV9K+hZoqHaQO5c3lHsqQtZG0BLyrjlAqMm/7JstdcywiO9BwuOLjz/R
vI3rI0Nh0hPTPoWh2h4ZiaM64K3EQ4whh7kdnoVpF2Ttl1PSCcZ1CQnxlyM4TBHR
g+f4zF67QkZ0F2pAIeN0Tv+qfhgDEWXl6dubJM5cYH4EM08QArJJ0R44y3GFvMPQ
A2PX1/l+8d990/UVPb+ZWs3i/9aP20R/gXybyTQDYUe3TmilwYOZwcNetRe4qc37
81gdsJSBV2mMcPOy4QTegVohoLs1IX6+wV1Sq3cRzw3CovtPJR68kz7YEJfsEQBO
FAoc20v4K1+8AVAFiNv2RK+O1HDpDtjNiJOa5LJNqeW0L7EfdzelrQAHLvNG88Ad
UYYFwo5VZXGk3k7u56hVVaDiaUqspnaxip7WUHmr9CvmLMpFa5T56yOPcHogfm2w
WT2+CvDZ++1h330a34SzxJNd91TwJvIMXuhN+G+x4EzJHthJ58dmuvUW+A84aIee
uLVR1q883QawzfrDLSKnv4gXHMn/Q8Iee5UfEc7DoQg7DgDAVgbFRhV8P8aZD4nd
VxnjirW9GGGiFaC8u4nZnYs/h5HFUicXY4cMNiBbJpAgYpD42f/JbCSlYCoAlYaM
VIZG3jBr5FfLjf5ewfTYlMD2jR4tQCovgRnEeBkFxgWJf2sFBTRH9BttVOgRGlMc
CGDWfwDjQDX4idGkrFBKUphK9ZORq9locJS4/X5WjPKNbX4NMPKFjeiYvs1saS1X
zXCk49EduKJoKnO1+ltOZMN8PrcM6CZFr8fmZgjXJ2mwDwd7fIjj2yfeH/aW+ruR
zJlrjrXWMMgV+3MLxhL3wJ+4H2qpON1aQDGl/Dstn4VDXTk+nrKcLBi+ur1kXlE+
Xa46BLY8HyILQHtLJU1hAbv9bJt/XnzyHJinmphDuQJCE9jRP+lRKl4nLIqJpT8G
PWx4jIobYXyInjQjnaFK3I+gdXftXVbK49I7DHnU/PiQA91KYx74woaE5XyRz5q8
EIi8jYQhFpXhBMKDJHykC8MTAxKPvr0CsnGwq8p3mbNtyWYf3liLYUEHC9tjgjrf
uhzqIlgz4j9CyVVBwWrOKiqH1YWLK3aXbxh0lUFtvDk+bBW+PmjzHmVcMCYxogFy
b387FjW1eyQ+gJ6oEbbNV3ylmUohfaVoNFAuwqeJENjoINDju2p0zQYRTbq2Zh17
OAze0AihABvCEKOUD+IhobFwijkEGc+EQeWxh+2dvSOebKqFufI9NZr4YERAr4th
pb9ss+yiAd3bbJroci9temc+gCALvJQhJtbOEr9H511CsYiv/Y8gshplvMnUwoqY
7RDnCODzHyyd3yFgELlmN/7Y54Y3MXBWj/gNJscIFhDKRhAcNToN5QI+ooqVYHKk
4kFkdFqWWw12vDeqVGqydMsAh1Hhps/ZiSWvwajPSM9MlOk1SE5zViDiiv0Yo10U
nJw49HK0n1LXcONrqW/ywOvhUrSmZS4O5M/jxfkA4AOKimrXMaOqufstBnzVlbHt
jtuYxh980LT4meF2ngYienG65iq+OSt7TPSXDMljkkbOGB4o5ra/RN9kZ7KiGgZA
PphR0e/EcUJxCoQeVuwE90lw6qCVFy3ItvNaJDLh7D3S61gkzaExZ7eRUy63wwLg
vzAz9k4CyCHQxnKpKNpzKTXYrGJfghEtsSNe87Xcga6jp6V3WAV1DP6OqpaDjGom
2P2ek+7hn4/u62tWWVYgGGlnyHRjFtwANow5GSHZAdtrNa90ATBPDj2g4evEs55j
v3z6ZVNDLxAYrPjP6LFEiWDg1ybG4z8EkK6nfuZialDNYlcEdV7d5qwiFTgVvK/T
h/NiO+EPmvk/d0C2TdKc/9+shlVpp5a1RYGYBBZzOQMcZwfmXDhR1KMgKWv2B3fM
hQH6O5p1ALLnL6KJe4ZNIAsYhq4Nu7KWhOFcwytX+8Ix6aTytt8NWYzCFAg7ryLo
wpIMVF7cj71uFmQ5eyJ29LNj7cTWZi1QE9s3q3HTwQU2egltyjzmCGWv567kjR7b
J4gfDG113stVmW6TskQmpdnbiomSxv97X91OJyyfQZWkO24bbL99hYb7Eyf5yFGM
vH/Ujr9ob6oKfM6W+VkemDJCYGpk+nZ2WmYuW+/wwKX5HNXOuZ83leX+sCuq0tjS
iWkiNyfaftkO8UGFSd+KMbwsK8VUiRKalAmYsg0NH3Zs+0XQPj5mpJqYyoa7K2ka
+gU2gly+5KMga3n1NWO98Y0CFBrAScX+RnvZo4DPZ3kWQSA/rygKOGTSXFkRmRw6
Kflmz+7a8BkwSVQzraiQ3LV/IpL7kYTgxaVrqim3cvKMcq2CFUkrS+dW71+Vvpsf
ZBFvjYAxrMOdERtUSjqVTneMKT/q0j21Rp/d+DZfGysWX8F+H6F2IT5QS4eZnwSV
4sjEEssQQWo8KFX93+g2qlmtAdcalN3H7UIITJbd2m+THaFcCcBfOJLJIKI8znbQ
YNMbnvwVW+f3ioB4br5ID9x8hJIabUPCexlevOgc//jcRmR6HJro1PQBZ753/avv
ZH9mVMXQJJJW3FrCfSYgUeWXo/0jXM2Ul+HJ7X9e7l4nP5Fz6on7q2fjoOWzcOCr
kGMcomBqb0syimWg2UGnAxMKOqp3QOUaGLySKgyYM5se2eAcIITt4BuFyxnVKH4Z
YfSO7j/2AcH2oddv1BBZWONtohm45tFQnfHatWMaUnxn/m6fKBy6pOT/HCY3c2Vq
7tvq1BOfuOSddmKMB/EElsM6fAKpUtoMKda5IbPVyZ+VBitk7Iku1lHmYqJfbWMM
G8X6C+v05ADK0muA12i3G19X39m7jZ4dRRPBZCqK6i66fX/jyXp2JrBur6Cdzm3G
rXDLtkFwAeZZrOsC9uOsaEYCl11lY44oA+c9lndnLF7xjTOQy27qeWOWtVEu7OQs
UliOHv3GYpYjwjc61ANehgEKCQTCfAdVtXhCtHFvWHWB7uSJv85lkw+Ky+ypi3oU
yW5Riqs/kDvInjjvLc8DOLE7qUEQceclElgRLdZ4hQn1LsWtaAvXML1ZrGXs6Aa1
ZObO2l/7VE/YHdOlVyJ2Ulrf8j7xaE3//Bs0tf3XaZyYLAhf8uvM7M7TU9KsGhSm
CAeC7pJXlhA4za93n7gK5QtOY+n/dBOQaVvyM5+LuupzkFY9jpCz1OCse+UTuIAq
56bC3cbHok+ElCA6JT1Uk9mPIYq4WBtxCFRsR5bzdbC7xnBHqVPp40fmOxQCp4Gp
8rGKNFLYkPIvERDVMWpq0OR5+6aVrFMi2LP/+FG5vFCqeczHrI/NNV56lh1ma0S/
bcT3SJu/5In+gFVDSUhf2OMeMHxfkgcb4hfxLAGitBf8hvoxt7z/6qskWp34FdtK
8ZGz1bInCV3akXdgeBTIKqlXKTnCaNROEpdoo9Heum7hMv5U3N7MDTU7qHyT4GRP
H6HMTEyGZpY/U8W2YnzVFGUwu7Z6lAoQuB+jjx+TNaFIb+UNNLvabWSjit9Ffcd1
5Wbfl+/8h5cCwEpsbO0Z0ZnKjYGJanPyaFIOwrKy6XQ+PYCvJs0hCvO9nQNHHCEu
PMt6a+0Lud+YHYLyMZ+ZQchFmPYpF4jUSzLj6FFo3P3ogfnaoluGVRoYlPUghRWe
Y/g1yndB03aSS46IJr8efn0MlgkCNLgOcncTE80zhwRp2cigDCF83LLQjQ9cf+Qu
oc6xH13H0YAAJq+fXWc2UyrL/1NmFcOEV9Dd9W5evAWjG+/ErcA4ta3YQ+q5KhH5
gy82sAwQ+ZLXkJhq5z8IvKeE1gIWL80h54xkCKHrDBtGoBBaAYLl8e8uAKRHs5ee
ue4iA2HnJAAWsqy+dDuTXOVmmGnzCyn9xpW0pNDR+0fx3o4PcGUcUy4ccNW2mLuG
3JV8hUQy0Yo438H4Lj//sIBCKanVvsDoCPjTko0iDDZI2rP/k4PwZuZ5+h4liJuE
N9oHafMj27eBh1TeS0vBMDTpr3kZK9lGVblOwknvoy8XbFZ8bZHzvpxc7JfLWUSk
n9fRgvuz+DS68nx+Tr6dApELpjC8OrLEgCwC5lzkk/ZQSEQTRYv68/2JI8TTEaxP
WcYrB4nUcjHH7np0DO25SgiiaQqSTUKXqN9Dlxal1/vPPlDU+CZMtRB5RR7S3zQm
+2LHtrSA3FDl6I4tEfbQdUDQlNixSuxmVskaPgBIc1Nd43WbaIDbj3S94FJ5Bcc1
FTvQGahw5wJaNQRwbcjYuA5F2du5bKDwK30eSfgQFEXAfJfLHP0/uoOOpUsyC3no
CE6Wbx+aHG3GFFxkCAZWFHEz6/ic18I4If4NMMQ5xs1EivYqMpK/fh7AwRpQvuiX
K0KVKB+J8oYOubWHPNsJkU3IKxC7Va3Mg7umFAV5vbsocuBW5ehNfBrWEKIEvHGV
tjcLmnNaLrNFgnPqfu4O/tQ4flHylMrT3+kE0Q2h9SYAOzpNDXOcfgh9NIJYR77Q
FYqzy45IcOsTfBhuOkcWIUOu6+H2ePXuDOI1YG5c79wCgGrD5BXdv6QRa+C5JdoI
cWA1Q548B1s2ldXLatXhWzUslGVlpVj5oISVWY3BrsWjCc2lBADR0G7fLuvYQisQ
TZt2rrqmTRsMVcWn7xdAS0jJpF6AOnPJP4XSbQ/TUHzsqj0Okpa09RBea8laPHnP
XdcMsrwVaQ/MVXQGLQEzw5riZjooU16hLpe8tGw54HVwfw5no7ChdD1Bo678Vgvk
gZO5Hqtw9gV53qQ7HeH+fnWRwaESrhSnhVuxeHCdkYXpDy6fVFDu6H+oWfQrirlK
O85QE6iH9rADPgDprFTn8y0Io/GpuOu1DcBbJaTsROM+pyyO9hr923Jar5c4DLpq
p+PYo3LLiP8wN+1snl8Z11tdXeGU1Kkr9aWoKzJzaVf0uHB+wdO/S/lUyFIKr099
9P7igQEwt8/P6hUE99T9zxErMRPf3pudYCV2Mhd9S+79thViWSjHNKhkYPWuyvvA
AlV29hw4vH2Gw/9TzBFZ6FsrP1XLXoQXVc9VVxZ9cQFNjeJd9xuNcj5ZRCEgHCvT
7qdb8B/E6iaaSTA8vcLP2Dh8ft4CelMveZBq1420gL10Ndv2A4DgquC+qKLNmowa
jUfj2S+nS18rlPdqwf5JZfhFoBHSDTDX/hiwh5J3f4VcmXUkrProY+jjMg4F/TZR
FNcqqN3iFRCqz+yxmh0/wPWfrhmaPwnD8JEzSPcLXpWDZWdYQH2KFQp6o8uT7LYY
uZAT7qq9Z9XXgO3qwsq9tPQQJAZzznYvTrLoA5DtnF//0HsmALZ1tccfoWKMq/l5
eD2+l1KrZb4LMEn5aY3H44RoxIu58KN/h6kHsf75UyIkibG/9WsUyGHq9fTlbERP
L94FHnGzQHUnOhZteZ6Iti6Y1FiXm60QWr4ibNDILlnHgQpFdmjwSoUye5pl76qi
GKcii6r1HwtD8RBTN98dSsOzafJvY1k1yezg5JMuUx/6dm3cBaH9udWNU4u14RKE
pCJsCQk8c0XSAnn6GEXPH1T2Swzy28LkYYSxSdSeistcd+U1O/Mzg3rE47tBtpZO
7s3K4f+3k96vXWhfu+bT+qE1sbIvcd/ki2DQCTBhqZ49mNfryCberxQ/XcJA05YC
3KzqXkjG26QAb/P5dg0wj0FrU/fqDc8khoCZGwS6NkanXlS2uueSDdicxajy2zQf
2Stwwg/Uv6Mc4lalz9SCgHjUqzaLM4rEiS+5frDujLKnfeAmw9zxvfuxRsIuswNo
QMiGoDrQc8jlBk7DtSX7pNlx0l15nfNo7qiEROPoksRGLUQubtH8ubJY8dik8seE
+SfEf8Rj24JVimoFgtcd+XLqxc443az/JvR0B32T8QH42uuiOfp5aPJVTIR3MhVY
Qp48mSVwj7cWYC2eTosFRMXjAjFcXrE73bf4v3Br9uN7RvPbEEWzNgWnzhA33a+/
KfVEFoeL6XK/S2YlU4GkXdFRQyQioc35W5+xBGRabMaZRp/MXdvZUzz80Bg6yLV6
6gLcEWZywCkuZO6f5uHpZ0NQhYBHZoF3iTtli3MBSE4VmH8ZhgzsZ67CvN2d1XEU
DrE2QqNFaeCDMt1ZIOoXLP5U7eivrjB8O7E3J03UAoXT2jApx3s6Kz/b/pptoOB6
Sg2V4mV2JDyFJuxwXbcW7sFvd58niWr64G36NazvqBuFvjaOK3MrpGK/ceDZYAQS
h5FJwGvB9dcMiSdOyzpsYKlzM1wAOf0lw9j2A0xdVJ5cUmNIqpqUpvlL+DdjB9+T
/IURWUkzpTPQweZejgd4k227hHNmLTFRObs3Csp/QpnrWKCaMjEt1O1ZB+Z+lQTz
mENxV08zFPN6ZE2B8OxAN4l2NypE27ITjY+yAnrX9dah+ZKaTu3ISmH9TLyvYDaM
vDhiX+CrELvfUYPEX6uShCd08xOwAscpM5+NHCJwoLCqWW2RT2sCD6RnAsIb1DLW
xx4u/KORGD0ew2YA2GcXzdoBIGv6pm1mwYqWlemb1xS8J2RKPjiCOfaRE4RA3IpN
LrrZ7o9hb3ukfz4RgchpJSC24MnteF7CHP4aDfsNF9/WUUPh4cEcULf4XJZtxrqf
kiGpr7M44WU1p2jwZRnptrpyB4MBvSbletakJn8O0SJv/zr5lgaa8B61fzSi7SYw
7jdzmp/yANA1ZsNy14RLkH8yYIYJ9VN21Lj4u6Y5LttBiLlEpKa63GqEpr2/U7Sy
XXxVoA3frrH38oxMVbwISIdJP0EN5qtqmoQ5+jKSgIPTPAVfXP02tVlmbxX61R5Y
8c3cGBHa0n23zquGnDNfGE8qjPQ+fGMvsNYZyBH4CtCWGDLhNs53sXcPWD2bbMfX
YwbbQUobXD+34Tz6j5QjunD5syLBSvz3EF44lN6FSlZtSUO8cVNLMfEi31ZvSB1Z
IQiG1y6i0j6lUxVcbFXL5ieNIcdFVpBhxi2QN7mHBXLDgj03QspHuPAtvWk3BKcQ
F7bP3L9sPnRPkg3PvNU5+J82uiFzh4cej4SjRnZvyCIMnRhGb8zVSO5EJkL120ET
8riifPae/65Ex8gxKossox+YOF/xpp9ZDoF2aixVkjcAo7M1jkXr2iE+0D6OCVhj
PAf4tgNaHlLLMNOrG6544Czd3DiOhH/DlI75iuGu0yTIrrdvrNjiqXy1hegX7rGc
85n6guQ7js3BNXZ5NUMKos2gSJqnZUusB5vv5CHslStVliQtagHuYBVxA+XCp29X
s628eT84fw9S+HmZuDHkihCnF4SwUY9P/D6GI9bFVvyCgusvXxJyvC2lcz84qsfm
6SBkEbb13rv00dXz9DtKAiEfbmNywBMPulYk7lmgWaJGxg/c+BPjs3quAlOqyYUt
jmN13wXffX72ZFKMgivCj7yxmipc2F3YNOAFsk+SNb2voNm6h0vhzTIZ0uEMOMpu
vQPEOwrkx3iVKrhqm485Gu7z/l46LMsCZ4GXSCzpgThLq34ezxBgnfWtOCy1i+9c
4ks27XpZU8tiQAWRZ+UKe3wiJXzKiC70VBG2Y4BSM10bHrD/mtkBti2jzqRts1qr
fVm1cpQnh3eI9X4UuLkl1xxe6awN96JNUE0m4xMWq9lz66K7j9zqy/gW57ES0p1D
uRiDtL/qjmqDhBjCAC2Otrlrf8pvJB3odaz2QR+dZ770d0lqBF7ceI+UL3+GqWHG
aq+cX1NkrPdfELC0cT573MqOCP5aQ7TJLcTwvhqiuyep9Vn9kSv7OeenI1zC9urm
Jm2cplHel0GVCpKBRqUWyYAKy1eJEvHvAaqei/iVGPCPywXKHgkLXJ2N6N0yDl5u
AKFnYJ6R94ZPBVklQ7MtKqzpX5u5If+tmQbxEHVaIfBoGaN/743DbCTuooYWLJsY
4I84azUwD6hrQJnjonqBTfjHb3qXZkYrbqwkmNge14a+6Ku4OJ6kjCsI/0ll5FdB
lE64GiTi+a/pzi0rZrUEARh5tklSM/alxusjAWpKYadjH3CmhQTt4yxoI2z3ALsS
Z4Gkz09qjx/v9ZQguu+yN9nuCMtWG1AOu73S1E9QmrkccyuctGLvCtkdFrGAgjSE
OjaTwjzhYwWO6kDzuF1s8/UGhkG2fs6Kr/825OPg44lWqX+OrZ0jUcCNCEdKlSdi
ftKavFX3mEJnSazn2n7qJPfc/JStnpDB+ZHriOdn+N60X2uTE8wFCKQXNZK0G7nI
c+9TKKqcY3VRma+inmeFO/4MSmFxhdvkDbNtQaynN6eUSIfy1KT4Xf1GEz/ymRrU
Mie4XkjK/L28DouECmfQY0idGJnij1HLifLpIleORXebRYLvek1bBzI2p20WHvam
wkpi1gUn1GQFSRMFaEHxtQivEMvpENNvwQoSjO/w5gIO2NDnOS5ccJuPkph5WV49
BynwruljeaMIWTqrXNnlJPPG1MapeRPtK+FYdEZSLnOzZ+KQfxe0mx54khszWxH3
Kclz6lD7NglHOXgtTfGU3lAdECNaKZc4BTuARfzVhFvQ00fzwsPCaraTu9vvFy4g
OwatYC/YshwoAbl91tdnVYXfRyfm1ABVPDq86lT80N6Y7BXQ8j5M1SnelSlRcFZL
zB6A3UnoA2sC+F5GdVGfMZ0OfJmkKywSeeO3m74t7nEs5x4+lnBX/pyMb9pPolBZ
kesEK4OYy7u0bg4EyqdIoUqxTMZ4vYgokwR3hVtgZDDIZjXSqLS7cVA4/IyODhP/
vrmr0qzJ1PARvNCFbb+OWyckKi53bTuczIFuBQvmE5OKyrbmqD8VeJf3Z6c5lFAk
Z1/fJ2v59uKOFof0Ss9KpDHycH6p09W7PoV4Sem15EwaT5ROtnG5aeL0tuxTgCeI
tl9zld3T6mnTs5BqcQpQvtwRbde7LN8kaG08oNDCcO4YzYm582C2BjnuVoTl2d0j
bMAKSDHpxBkNMQvpORCRi033Hcr0M9lyVXZ7icqcvea0hzAFRASNp9BP4qGU+9wT
p1ux8OnjSJEpJrcMtJ1Kt2Qpsr7kZ1AVx9IhQMJPRRlYiHo3iuIulR3dfUipMfrd
v0MK7EfutKAIhMDRAasK1ohpiYtc3a16KefMIB2v8P1IMyJx9kv5lXjW9rzHNDnp
DuhORfSYEnNNa0zG58o0oYfOobzqh5azeiTs9F8Lifp0CPMWQBV0kSZFcy+8OEHU
bb6E1fQoz9/lfPuqVxXPAUaqVqbZTzUnDYSwgx07XQf1WkIiwlvcnW8Y6zCqMP9X
F9h7xjt+ez64U8YJRrFlEQJAnU/2UQyRPodV6BGjq96dSGccQQnmsCGSokQGVE28
ziA6AfbNeWFUEK2TjKYks7tZDs9gv+xN05aszMwJdU015tfs0LwEE7GULSyQJCyU
Cl2Uc5/NJV3LYJJH29VwrDb+1T4o4BT7qnA0vCgVFEmNQ3Kvoul3ZQpFTCoNiL6e
ktEotcKN/+7dYMGwa+sVFxkgvWzURCrIJAdOKUaAic8+N3aKpj2MFMetp2473RA9
4FuVPLeUX8rD1iTeOYG4VE7NQbVgwH5jBaUNwMi0i4RVM1ZP8O9UkgfDokIHb5br
m6TlLd1z/h+vCy6/7aIlRuogROhfpGlWHHTXJakd+DSd6elrg553/PckbyqTkjh7
uH00LcA/r0jeMuNFCg0S5nmILHzDBH6TUVI7Lngrpe9oOcfMs5b7zquutWi32y+v
DY7pifHUCobS/kLHzMx8kNq/UwTG/8cO5nWlnOtTbbnyHasyOHB8ZtfHJYeKxSPz
bF80KcPJ8W+p+JG/OZSTd0lXaCYZ95RS6UyH7BleveptZAT5lXAgaW4va3r+uneD
ziBLbEF+chlkz9HMFaEnNrZVYoun1Lus1xBu9zDzZdGdrj55k2dpeRYBSCnXUimi
C4HKKKqKwCGlVsX50EdYc9yDYiBsWLpkKi0E+XJDFZGOjB322OY1MuteqSSyg1YX
yjVfCWdDiDENI6mEZ1Sc2zX/Pz45huNl/ITnouZ2mGkyEQRhAI2tT8SsJkfwhZcc
2ZK+ZNWO/HodKMe5JiTqKHQdTP16H+w3vKCVmvV9Lr6rTTEhGab9JeihMKfGqJBs
6Z2YVPXJGgQbbiR1pKOFKQI9FnwR1cYzrnmZ4Rwbwt0flJe/e0fTz793IpHEursc
U/QZviSo91DYlDOIy8A/2Nql/RQNkcCw4gzqE3MRoJZSvz0yvss8p6MVwSFPIyR0
IPoZTK2u7+M9HTON85iQWvzQ9AIbUriOwPV/O2eydkHj2DJRpUmQ6vNUnxyw+xnb
Wz/04latwquutiCg0yeqDEdDOJG/QbAWqdBMkcXi8waWN/31abumWYWarHKDtDsd
`pragma protect end_protected
