// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cyRv8JRFIS8YHu534yLdkJ7MFgeaTGo9qECPobjuu9+YBwr4KDn1VF43Vuytvjy1
901vlwB9q4/r6+RE7c7rS8K3SRg7dDJ6uK9hluybwa7IUaMA1f2B0LlcrLwQqFJE
pvEK6c7IFDRqjP4rgk2hnnNdlez4u//GQSkANwlbmag=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2368)
e9WTVYLtqDzzz6UZuB+zxrsXkMiUTn6uK/NOvg1/wbAJQtJZL1gEzKMHb5nfBPvU
3OiBnWmNLULHo/3nZioSYDYsRn76j7OIlGKahQD8N7G5U3cSIslKZqPg/SrNIx4M
xaKk5EwFbKSFcxABrZ1id+jv48iajYkB5sb9a0C7eqi2MFJtjaMk1WxSfAvRPmiA
Dvam3Lv0bI93f7jXuShvNfIZHG79oK4OA515ofBXdLUlOyFTEvMPkmmdSbm0QD3O
RgD1KUD5vjYotlaL58uHFORjp1o/X+Li3sPjwtSflyLqZbR9OaoEKr8/CUVYwmhR
6oyEP4DEVjJeiokGZlYKrZHfj91JT9n233MTuG0O03/jRlwy1+fLnRV/GihDPGvL
rXzKxEDyUxz238qHtnSdCVrzg68iJBcbfRqF0ZUAv9FnkorshGyjrb3lqI+F6skk
v3xA6CSRl8sRzbP6xDlj4FE+MBRjpZlImhURUcmeKY1+sOBCs3Lg4Pig+1aILiEB
J6V0TzUomTCNQ2pUVnswZ7yee/zvsGH4Hs89o3GpAQ6ATl1QCsuVsJF26GxeeYFL
xvjbzksH+sOUQmgtxQzrrnnJN/15UOIfR3XKEaHKxRsriaaHtl52ENmmU7xErwjd
+MmzoDBqGtDQZiTblhq5btABcqDyee05Ct4SslUneH9Bxngcaa/TBopiI/clXFJu
7vAFHwMRZQ9EH3bZLkJoZSa2CsdtIlQIzMHz/iEGVMl8/maWIDayMp+BwIT4w/ok
7LoZ52gBZ4KZiGw4cBv4DxtbX2xFSuGSEDpH79PIZ3bCBuLVypEsvhKv7W+QORWv
+L7udFk/uqgp3dpF7TwKCyEr8/I96r9m3CEGvP+hMkMIkfMowewhylGKzhON+ASJ
H+3i6eubPCdEcg8r1My6a7iKTd9obsdNzFw/ku2e15CU4YFYM43eJ9O/clpOWa3Q
2PmPDEFHWmPlX2VCGi65pOo4cNpo+xMJMtlOFj+sMcP71qiLjYjfPY0bNMi1N+es
C349WdLHkphws2aP9NP4/hXi2w9n82KV5eoBbh47suaVKrfySu0WL/ttAyGghAW+
AsJDL7kO0ckhS9h26NRLLLxV44lhIp2uY6pAeTzgAWdUfd4ZuTU4FJOkZcbOmIdS
6WRliMuMW3e8AlwB9BNhCmO4Z1NeQWr6ZiUPeHXQrguXfRGAEG5MWKO6jMvRHrLY
CZVwSQyqIQb/8JNdBEgmY/CSS/53xS2XGQAi1U7EvT/Td9dg4RFddqC5QqHzQzSW
vOzY2ZBsKsY2/rdcfIVG+11CaJ4TFL30kwP4nRQ/SiV6v9rb8MF6YSXf8AkUFpec
tN/Ylf5VHw6QYXvPP7Ayj2UjhgKPVvKcMZs3RAXevQMmi4mdeCUuyAwxbNZfCHk6
qwlBMjDrBPJ1N5N34ojn0niUW5gSlMJSC3SYfEpH7zOAFAgV3j5hcHJFGuUu5pFt
vLszhxbNqSp1qTlANAdQjhwIG5K8e4IylkZikbtIhq+i51aVrmYBcTgGXeNrd8Qh
qTJ6IXpc8C94tV6/hPz2dttOTMTQQJKgsq7xfMUr0jxItyse4qHtMMjTBDYyQ+Em
DVv6gW4tZwC8t3+Ss+exJNql0j9PUtVI+6FU+pVBIS0PpkEQrwgPwCxZFP12kUmA
ApdXww9PrK00CxjpugihcbyBd5aK81kBVKruwvqXx3cO/HxH3r2MusHH0OrijB0y
TLyUk+TrJ4ikn56+3UbY8PfgeQkS+GOvDEbOv5riKj9ND7r0vpZa8ehuh5Zhw0uC
/yJbjdXlLn4FpfNnCS8TbNNzowFfVCOcIvUCBlv/eow5dqYmIakvn1nfW7j40XFf
9mCAMYxEXpUX/O1Qs8imaxpw7eAH0ZgQNtmNvjnP3b38o7Hl0jqR7zm8P8unly6a
XdRPLmSGlqCMqBJ8+1Rjx19FPP/ekIaj/c8/iGk6Kc+NFJjFxyoLyeIvR06k09AI
i+TQaIuiclHVzNIKaztFsHkKWczK8q0usyNLtSjqvqFq3CRxv4UMdq80n22+SjNr
6VpXWpMtAKMqSwwceHA3gHQqCBCqPC9Z7+qOwInoHzWjrE3jfCsFPg9jGhjOx8lD
1qdHn9H1q41pINqwZhZi7jAhi4Q5s3mstRa3SLE29uqzU80yhaEEzs+8jzDzRunD
IyNipZ3BZaezl74cYleKhPsAXzxe7EEN9/VBAu1GY29OnmzPWp9TNiKqZ9SN9moP
lbhD9NY0iIdGW+bIghoWYhibf45ExC8BOMUBVCJMWRrXYn29X4fz9IKvDRmi48w+
XGm+7e3bwmR04qTceA/O5poZm3o4l/2iBsgtJpojTabv8hKatBmpHslqxB0D4p3v
fecUbQ1I0wmD4BOcJA4FljsYV8NP0VMXXABKUYUFwXyBcJ2CvcAGJMgonMJKfhqu
OihQX4XKY27DJwrrIBJkhPBZrlB1gkekTEu8rFqKN0EfU8jjZafKpUxRjNLEQyfj
xZ8R4S8kZljYK2WabmK1ZXP8MPUKX0xM+wDQ7gy3sqPIO79OIChh2f9Eyced5GA6
jJePR8vhzobpv6mNqiBPaurGS3dRaqXqpm2xrdqpUgHEoicGhIM6d31hH7M+FETR
8HzXoRYDDyImbMXMS2czBACf6+FXu2s3AivdEvatx/0CQuD7ipT7PnybMkw6gYi4
SyxiLMOp+QgU4iFWWPeSsPi6Gq0DPUyd5zl+Gpakwz/WDnrOsDhNp2ySF5+VeQFM
mY9hiL65cJuz+ZH3FZOGPVnZN1TIlkYlbpnswmSdeOXOJkwK9uYpYM8OAIMySCe/
sb0aYWX7jsssztpI3gYg+KZc5Gp10/nVnlVVa7va8CcKVjstEvUpVVxmPNZKZHwV
CUG42V4klEfvUKZARG1JirXbUhzqRZy+zE7LdTIZhZKNXwnYM+YcofkTPBpSm8Rh
+XyHaRxjbuYRvw6qY5QKNfoliu6+OYrat61kDhmy9JEiNcrp81LgsivJC3NcnhRD
1EftpHS1IAbyyHzBffZB15eMPVQPCMvo2EIOuCkI6W/Jlr5inqDYT00Obnih2hhL
a3TuvjE7cJ0u82qK6g7EdUPCOY7als+92qC6gqhUKauofD7cG5luaKAi1jGo2qMm
Ufa33xSlKyFXTgmObQcw9A==
`pragma protect end_protected
